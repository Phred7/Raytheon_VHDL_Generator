library IEEE;
    use IEEE.std_logic_1164.all;
    use IEEE.numeric_std.all;
    package lowlife_package is
    constant FORMAT_2 : integer := 15;
    constant JMP1 : integer := 0;
    constant JMP2 : integer := 1;
    constant MOV : integer := 2;
    constant OFFSET : integer := -2;
    end lowlife_package;
