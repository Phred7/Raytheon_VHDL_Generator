library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;


entity highroller_memory is
    port ( clk	: in	std_logic;
         MAB		: in	std_logic_vector(15 downto 0);
         MDB_in  	: out	std_logic_vector(15 downto 0);
         MDB_out  	: in	std_logic_vector(15 downto 0);
         write	    : in	std_logic);
end entity;

architecture highroller_memory_arch of highroller_memory is

type rom_type is array (32768 to 65535) of std_logic_vector(7 downto 0);  -- this is MAB: x8000 to xFFFF
    
constant ROM : rom_type :=(						   55896 => x"B2",		-- 00da58: B240             MOV.W   #0x5a80,&WDTCTL_L
						   55897 => x"60",
						   55898 => x"80",		-- 00da5a: 805A            
						   55899 => x"5A",
						   55900 => x"CC",		-- 00da5c: CC01            
						   55901 => x"01",
						   55902 => x"91",		-- 00da5e: 9142             MOV.W   &$P$T0$1,0x0002(SP)
						   55903 => x"62",
						   55904 => x"3E",		-- 00da60: 3E9A            
						   55905 => x"9A",
						   55906 => x"02",		-- 00da62: 0200            
						   55907 => x"00",
						   55908 => x"91",		-- 00da64: 9142             MOV.W   &0x9a40,0x0004(SP)
						   55909 => x"62",
						   55910 => x"40",		-- 00da66: 409A            
						   55911 => x"9A",
						   55912 => x"04",		-- 00da68: 0400            
						   55913 => x"00",
						   55914 => x"91",		-- 00da6a: 9142             MOV.W   &0x9a42,0x0006(SP)
						   55915 => x"62",
						   55916 => x"42",		-- 00da6c: 429A            
						   55917 => x"9A",
						   55918 => x"06",		-- 00da6e: 0600            
						   55919 => x"00",
						   55920 => x"91",		-- 00da70: 9142             MOV.W   &0x9a44,0x0008(SP)
						   55921 => x"62",
						   55922 => x"44",		-- 00da72: 449A            
						   55923 => x"9A",
						   55924 => x"08",		-- 00da74: 0800            
						   55925 => x"00",
						   55926 => x"81",		-- 00da76: 8143             CLR.W   0x000a(SP)
						   55927 => x"63",
						   55928 => x"0A",		-- 00da78: 0A00            
						   55929 => x"00",
						   55930 => x"81",		-- 00da7a: 8193             TST.W   0x000a(SP)
						   55931 => x"B3",
						   55932 => x"0A",		-- 00da7c: 0A00            
						   55933 => x"00",
						   55934 => x"06",		-- 00da7e: 0620             JNE     ($C$L1)
						   55935 => x"40",
						   55936 => x"B1",		-- 00da80: B140             MOV.W   #0x8514,0x0000(SP)
						   55937 => x"60",
						   55938 => x"14",		-- 00da82: 1485            
						   55939 => x"85",
						   55940 => x"00",		-- 00da84: 0000            
						   55941 => x"00",
						   55942 => x"B0",		-- 00da86: B012             CALL    #printf
						   55943 => x"32",
						   55944 => x"EE",		-- 00da88: EEDC            
						   55945 => x"DC",
						   55946 => x"05",		-- 00da8a: 053C             JMP     ($C$L2)
						   55947 => x"5C",
						   55948 => x"B1",		-- 00da8c: B140             MOV.W   #0x8514,0x0000(SP)
						   55949 => x"60",
						   55950 => x"14",		-- 00da8e: 1485            
						   55951 => x"85",
						   55952 => x"00",		-- 00da90: 0000            
						   55953 => x"00",
						   55954 => x"B0",		-- 00da92: B012             CALL    #printf
						   55955 => x"32",
						   55956 => x"EE",		-- 00da94: EEDC            
						   55957 => x"DC",
						   55958 => x"0C",		-- 00da96: 0C43             CLR.W   R12
						   55959 => x"63",
						   55960 => x"31",		-- 00da98: 3150             ADD.W   #0x000c,SP
						   55961 => x"70",
						   55962 => x"0C",		-- 00da9a: 0C00            
						   55963 => x"00",
						   55964 => x"30",		-- 00da9c: 3041             RET     
						   55965 => x"61",
						   -- Begin: __mspabi_srlll
						   55966 => x"07",		-- 00da9e: 0712             PUSH    R7
						   55967 => x"32",
						   55968 => x"07",		-- 00daa0: 074C             MOV.W   R12,R7
						   55969 => x"6C",
						   55970 => x"0D",		-- 00daa2: 0D49             MOV.W   R9,R13
						   55971 => x"69",
						   55972 => x"0E",		-- 00daa4: 0E4A             MOV.W   R10,R14
						   55973 => x"6A",
						   55974 => x"0F",		-- 00daa6: 0F4B             MOV.W   R11,R15
						   55975 => x"6B",
						   55976 => x"37",		-- 00daa8: 3790             CMP.W   #0x0011,R7
						   55977 => x"B0",
						   55978 => x"11",		-- 00daaa: 1100            
						   55979 => x"00",
						   55980 => x"0E",		-- 00daac: 0E38             JL      ($C$L2)
						   55981 => x"58",
						   55982 => x"0B",		-- 00daae: 0B47             MOV.W   R7,R11
						   55983 => x"67",
						   55984 => x"1B",		-- 00dab0: 1B83             DEC.W   R11
						   55985 => x"A3",
						   55986 => x"0C",		-- 00dab2: 0C4B             MOV.W   R11,R12
						   55987 => x"6B",
						   55988 => x"B0",		-- 00dab4: B012             CALL    #__mspabi_srai_4
						   55989 => x"32",
						   55990 => x"6A",		-- 00dab6: 6ADE            
						   55991 => x"DE",
						   55992 => x"3B",		-- 00dab8: 3BF0             AND.W   #0xfff0,R11
						   55993 => x"10",
						   55994 => x"F0",		-- 00daba: F0FF            
						   55995 => x"FF",
						   55996 => x"07",		-- 00dabc: 078B             SUB.W   R11,R7
						   55997 => x"AB",
						   55998 => x"08",		-- 00dabe: 084D             MOV.W   R13,R8
						   55999 => x"6D",
						   56000 => x"0D",		-- 00dac0: 0D4E             MOV.W   R14,R13
						   56001 => x"6E",
						   56002 => x"0E",		-- 00dac2: 0E4F             MOV.W   R15,R14
						   56003 => x"6F",
						   56004 => x"0F",		-- 00dac4: 0F43             CLR.W   R15
						   56005 => x"63",
						   56006 => x"1C",		-- 00dac6: 1C83             DEC.W   R12
						   56007 => x"A3",
						   56008 => x"FA",		-- 00dac8: FA23             JNE     ($C$L1)
						   56009 => x"43",
						   56010 => x"17",		-- 00daca: 1793             CMP.W   #1,R7
						   56011 => x"B3",
						   56012 => x"08",		-- 00dacc: 0838             JL      ($C$L4)
						   56013 => x"58",
						   56014 => x"0C",		-- 00dace: 0C47             MOV.W   R7,R12
						   56015 => x"67",
						   56016 => x"12",		-- 00dad0: 12C3             CLRC    
						   56017 => x"E3",
						   56018 => x"0F",		-- 00dad2: 0F10             RRC     R15
						   56019 => x"30",
						   56020 => x"0E",		-- 00dad4: 0E10             RRC     R14
						   56021 => x"30",
						   56022 => x"0D",		-- 00dad6: 0D10             RRC     R13
						   56023 => x"30",
						   56024 => x"08",		-- 00dad8: 0810             RRC     R8
						   56025 => x"30",
						   56026 => x"1C",		-- 00dada: 1C83             DEC.W   R12
						   56027 => x"A3",
						   56028 => x"F9",		-- 00dadc: F923             JNE     ($C$L3)
						   56029 => x"43",
						   56030 => x"0C",		-- 00dade: 0C48             MOV.W   R8,R12
						   56031 => x"68",
						   56032 => x"37",		-- 00dae0: 3741             POP.W   R7
						   56033 => x"61",
						   56034 => x"30",		-- 00dae2: 3041             RET     
						   56035 => x"61",
						   -- Begin: HOSTclose
						   56036 => x"0A",		-- 00dae4: 0A12             PUSH    R10
						   56037 => x"32",
						   56038 => x"0A",		-- 00dae6: 0A4C             MOV.W   R12,R10
						   56039 => x"6C",
						   56040 => x"92",		-- 00dae8: 9212             CALL    &_lock
						   56041 => x"32",
						   56042 => x"F2",		-- 00daea: F220            
						   56043 => x"20",
						   56044 => x"C2",		-- 00daec: C24A             MOV.B   R10,&parmbuf
						   56045 => x"6A",
						   56046 => x"9E",		-- 00daee: 9E21            
						   56047 => x"21",
						   56048 => x"8A",		-- 00daf0: 8A10             SWPB    R10
						   56049 => x"30",
						   56050 => x"8A",		-- 00daf2: 8A11             SXT     R10
						   56051 => x"31",
						   56052 => x"C2",		-- 00daf4: C24A             MOV.B   R10,&0x219f
						   56053 => x"6A",
						   56054 => x"9F",		-- 00daf6: 9F21            
						   56055 => x"21",
						   56056 => x"7C",		-- 00daf8: 7C40             MOV.B   #0x00f1,R12
						   56057 => x"60",
						   56058 => x"F1",		-- 00dafa: F100            
						   56059 => x"00",
						   56060 => x"3D",		-- 00dafc: 3D40             MOV.W   #0x219e,R13
						   56061 => x"60",
						   56062 => x"9E",		-- 00dafe: 9E21            
						   56063 => x"21",
						   56064 => x"0E",		-- 00db00: 0E43             CLR.W   R14
						   56065 => x"63",
						   56066 => x"0F",		-- 00db02: 0F43             CLR.W   R15
						   56067 => x"63",
						   56068 => x"B0",		-- 00db04: B012             CALL    #__TI_writemsg
						   56069 => x"32",
						   56070 => x"92",		-- 00db06: 92DD            
						   56071 => x"DD",
						   56072 => x"3C",		-- 00db08: 3C40             MOV.W   #0x219e,R12
						   56073 => x"60",
						   56074 => x"9E",		-- 00db0a: 9E21            
						   56075 => x"21",
						   56076 => x"0D",		-- 00db0c: 0D43             CLR.W   R13
						   56077 => x"63",
						   56078 => x"B0",		-- 00db0e: B012             CALL    #__TI_readmsg
						   56079 => x"32",
						   56080 => x"1C",		-- 00db10: 1CDE            
						   56081 => x"DE",
						   56082 => x"5F",		-- 00db12: 5F42             MOV.B   &parmbuf,R15
						   56083 => x"62",
						   56084 => x"9E",		-- 00db14: 9E21            
						   56085 => x"21",
						   56086 => x"5A",		-- 00db16: 5A42             MOV.B   &0x219f,R10
						   56087 => x"62",
						   56088 => x"9F",		-- 00db18: 9F21            
						   56089 => x"21",
						   56090 => x"8A",		-- 00db1a: 8A10             SWPB    R10
						   56091 => x"30",
						   56092 => x"0A",		-- 00db1c: 0A5F             ADD.W   R15,R10
						   56093 => x"7F",
						   56094 => x"92",		-- 00db1e: 9212             CALL    &_unlock
						   56095 => x"32",
						   56096 => x"F4",		-- 00db20: F420            
						   56097 => x"20",
						   56098 => x"0C",		-- 00db22: 0C4A             MOV.W   R10,R12
						   56099 => x"6A",
						   56100 => x"3A",		-- 00db24: 3A41             POP.W   R10
						   56101 => x"61",
						   56102 => x"30",		-- 00db26: 3041             RET     
						   56103 => x"61",
						   -- Begin: __mspabi_sllll
						   56104 => x"07",		-- 00db28: 0712             PUSH    R7
						   56105 => x"32",
						   56106 => x"07",		-- 00db2a: 074C             MOV.W   R12,R7
						   56107 => x"6C",
						   56108 => x"0D",		-- 00db2c: 0D49             MOV.W   R9,R13
						   56109 => x"69",
						   56110 => x"0E",		-- 00db2e: 0E4A             MOV.W   R10,R14
						   56111 => x"6A",
						   56112 => x"0F",		-- 00db30: 0F4B             MOV.W   R11,R15
						   56113 => x"6B",
						   56114 => x"37",		-- 00db32: 3790             CMP.W   #0x0011,R7
						   56115 => x"B0",
						   56116 => x"11",		-- 00db34: 1100            
						   56117 => x"00",
						   56118 => x"0E",		-- 00db36: 0E38             JL      ($C$L2)
						   56119 => x"58",
						   56120 => x"0F",		-- 00db38: 0F47             MOV.W   R7,R15
						   56121 => x"67",
						   56122 => x"1F",		-- 00db3a: 1F83             DEC.W   R15
						   56123 => x"A3",
						   56124 => x"0C",		-- 00db3c: 0C4F             MOV.W   R15,R12
						   56125 => x"6F",
						   56126 => x"B0",		-- 00db3e: B012             CALL    #__mspabi_srai_4
						   56127 => x"32",
						   56128 => x"6A",		-- 00db40: 6ADE            
						   56129 => x"DE",
						   56130 => x"3F",		-- 00db42: 3FF0             AND.W   #0xfff0,R15
						   56131 => x"10",
						   56132 => x"F0",		-- 00db44: F0FF            
						   56133 => x"FF",
						   56134 => x"07",		-- 00db46: 078F             SUB.W   R15,R7
						   56135 => x"AF",
						   56136 => x"0F",		-- 00db48: 0F4E             MOV.W   R14,R15
						   56137 => x"6E",
						   56138 => x"0E",		-- 00db4a: 0E4D             MOV.W   R13,R14
						   56139 => x"6D",
						   56140 => x"0D",		-- 00db4c: 0D48             MOV.W   R8,R13
						   56141 => x"68",
						   56142 => x"08",		-- 00db4e: 0843             CLR.W   R8
						   56143 => x"63",
						   56144 => x"1C",		-- 00db50: 1C83             DEC.W   R12
						   56145 => x"A3",
						   56146 => x"FA",		-- 00db52: FA23             JNE     ($C$L1)
						   56147 => x"43",
						   56148 => x"17",		-- 00db54: 1793             CMP.W   #1,R7
						   56149 => x"B3",
						   56150 => x"07",		-- 00db56: 0738             JL      ($C$L4)
						   56151 => x"58",
						   56152 => x"0C",		-- 00db58: 0C47             MOV.W   R7,R12
						   56153 => x"67",
						   56154 => x"08",		-- 00db5a: 0858             RLA.W   R8
						   56155 => x"78",
						   56156 => x"0D",		-- 00db5c: 0D6D             RLC.W   R13
						   56157 => x"8D",
						   56158 => x"0E",		-- 00db5e: 0E6E             RLC.W   R14
						   56159 => x"8E",
						   56160 => x"0F",		-- 00db60: 0F6F             RLC.W   R15
						   56161 => x"8F",
						   56162 => x"1C",		-- 00db62: 1C83             DEC.W   R12
						   56163 => x"A3",
						   56164 => x"FA",		-- 00db64: FA23             JNE     ($C$L3)
						   56165 => x"43",
						   56166 => x"0C",		-- 00db66: 0C48             MOV.W   R8,R12
						   56167 => x"68",
						   56168 => x"37",		-- 00db68: 3741             POP.W   R7
						   56169 => x"61",
						   56170 => x"30",		-- 00db6a: 3041             RET     
						   56171 => x"61",
						   -- Begin: exit
						   56172 => x"0A",		-- 00db6c: 0A12             PUSH    R10
						   56173 => x"32",
						   56174 => x"0A",		-- 00db6e: 0A4C             MOV.W   R12,R10
						   56175 => x"6C",
						   56176 => x"82",		-- 00db70: 8293             TST.W   &__TI_enable_exit_profile_output
						   56177 => x"B3",
						   56178 => x"FA",		-- 00db72: FA20            
						   56179 => x"20",
						   56180 => x"0A",		-- 00db74: 0A24             JEQ     ($C$L3)
						   56181 => x"44",
						   56182 => x"3E",		-- 00db76: 3E40             MOV.W   #0xffff,R14
						   56183 => x"60",
						   56184 => x"FF",		-- 00db78: FFFF            
						   56185 => x"FF",
						   56186 => x"3F",		-- 00db7a: 3F40             MOV.W   #0xffff,R15
						   56187 => x"60",
						   56188 => x"FF",		-- 00db7c: FFFF            
						   56189 => x"FF",
						   56190 => x"3F",		-- 00db7e: 3F93             CMP.W   #-1,R15
						   56191 => x"B3",
						   56192 => x"02",		-- 00db80: 0220             JNE     ($C$L2)
						   56193 => x"40",
						   56194 => x"3E",		-- 00db82: 3E93             CMP.W   #-1,R14
						   56195 => x"B3",
						   56196 => x"02",		-- 00db84: 0224             JEQ     ($C$L3)
						   56197 => x"44",
						   56198 => x"B0",		-- 00db86: B012             CALL    #0xffff
						   56199 => x"32",
						   56200 => x"FF",		-- 00db88: FFFF            
						   56201 => x"FF",
						   56202 => x"92",		-- 00db8a: 9212             CALL    &_lock
						   56203 => x"32",
						   56204 => x"F2",		-- 00db8c: F220            
						   56205 => x"20",
						   56206 => x"82",		-- 00db8e: 8293             TST.W   &__TI_dtors_ptr
						   56207 => x"B3",
						   56208 => x"F0",		-- 00db90: F020            
						   56209 => x"20",
						   56210 => x"03",		-- 00db92: 0324             JEQ     ($C$L4)
						   56211 => x"44",
						   56212 => x"0C",		-- 00db94: 0C4A             MOV.W   R10,R12
						   56213 => x"6A",
						   56214 => x"92",		-- 00db96: 9212             CALL    &__TI_dtors_ptr
						   56215 => x"32",
						   56216 => x"F0",		-- 00db98: F020            
						   56217 => x"20",
						   56218 => x"82",		-- 00db9a: 8293             TST.W   &__TI_cleanup_ptr
						   56219 => x"B3",
						   56220 => x"EE",		-- 00db9c: EE20            
						   56221 => x"20",
						   56222 => x"02",		-- 00db9e: 0224             JEQ     ($C$L5)
						   56223 => x"44",
						   56224 => x"92",		-- 00dba0: 9212             CALL    &__TI_cleanup_ptr
						   56225 => x"32",
						   56226 => x"EE",		-- 00dba2: EE20            
						   56227 => x"20",
						   56228 => x"92",		-- 00dba4: 9212             CALL    &_unlock
						   56229 => x"32",
						   56230 => x"F4",		-- 00dba6: F420            
						   56231 => x"20",
						   56232 => x"B0",		-- 00dba8: B012             CALL    #abort
						   56233 => x"32",
						   56234 => x"B8",		-- 00dbaa: B8E1            
						   56235 => x"E1",
						   56236 => x"3A",		-- 00dbac: 3A41             POP.W   R10
						   56237 => x"61",
						   56238 => x"30",		-- 00dbae: 3041             RET     
						   56239 => x"61",
						   -- Begin: __TI_auto_init_nobinit_nopinit
						   56240 => x"0A",		-- 00dbb0: 0A12             PUSH    R10
						   56241 => x"32",
						   56242 => x"09",		-- 00dbb2: 0912             PUSH    R9
						   56243 => x"32",
						   56244 => x"3F",		-- 00dbb4: 3F40             MOV.W   #0x8502,R15
						   56245 => x"60",
						   56246 => x"02",		-- 00dbb6: 0285            
						   56247 => x"85",
						   56248 => x"3F",		-- 00dbb8: 3F90             CMP.W   #0x8508,R15
						   56249 => x"B0",
						   56250 => x"08",		-- 00dbba: 0885            
						   56251 => x"85",
						   56252 => x"16",		-- 00dbbc: 1624             JEQ     ($C$L22)
						   56253 => x"44",
						   56254 => x"3F",		-- 00dbbe: 3F40             MOV.W   #0x850c,R15
						   56255 => x"60",
						   56256 => x"0C",		-- 00dbc0: 0C85            
						   56257 => x"85",
						   56258 => x"3F",		-- 00dbc2: 3F90             CMP.W   #0x8514,R15
						   56259 => x"B0",
						   56260 => x"14",		-- 00dbc4: 1485            
						   56261 => x"85",
						   56262 => x"11",		-- 00dbc6: 1124             JEQ     ($C$L22)
						   56263 => x"44",
						   56264 => x"3A",		-- 00dbc8: 3A40             MOV.W   #0x8514,R10
						   56265 => x"60",
						   56266 => x"14",		-- 00dbca: 1485            
						   56267 => x"85",
						   56268 => x"3A",		-- 00dbcc: 3A80             SUB.W   #0x850c,R10
						   56269 => x"A0",
						   56270 => x"0C",		-- 00dbce: 0C85            
						   56271 => x"85",
						   56272 => x"0A",		-- 00dbd0: 0A11             RRA     R10
						   56273 => x"31",
						   56274 => x"0A",		-- 00dbd2: 0A11             RRA     R10
						   56275 => x"31",
						   56276 => x"39",		-- 00dbd4: 3940             MOV.W   #0x850c,R9
						   56277 => x"60",
						   56278 => x"0C",		-- 00dbd6: 0C85            
						   56279 => x"85",
						   56280 => x"3C",		-- 00dbd8: 3C49             MOV.W   @R9+,R12
						   56281 => x"69",
						   56282 => x"7F",		-- 00dbda: 7F4C             MOV.B   @R12+,R15
						   56283 => x"6C",
						   56284 => x"0F",		-- 00dbdc: 0F5F             RLA.W   R15
						   56285 => x"7F",
						   56286 => x"1F",		-- 00dbde: 1F4F             MOV.W   0x8502(R15),R15
						   56287 => x"6F",
						   56288 => x"02",		-- 00dbe0: 0285            
						   56289 => x"85",
						   56290 => x"3D",		-- 00dbe2: 3D49             MOV.W   @R9+,R13
						   56291 => x"69",
						   56292 => x"8F",		-- 00dbe4: 8F12             CALL    R15
						   56293 => x"32",
						   56294 => x"1A",		-- 00dbe6: 1A83             DEC.W   R10
						   56295 => x"A3",
						   56296 => x"F7",		-- 00dbe8: F723             JNE     ($C$L21)
						   56297 => x"43",
						   56298 => x"B0",		-- 00dbea: B012             CALL    #_system_post_cinit
						   56299 => x"32",
						   56300 => x"C8",		-- 00dbec: C8E1            
						   56301 => x"E1",
						   56302 => x"30",		-- 00dbee: 3040             BR      #__mspabi_func_epilog_2
						   56303 => x"60",
						   56304 => x"64",		-- 00dbf0: 64E1            
						   56305 => x"E1",
						   -- Begin: HOSTunlink
						   56306 => x"0A",		-- 00dbf2: 0A12             PUSH    R10
						   56307 => x"32",
						   56308 => x"0A",		-- 00dbf4: 0A4C             MOV.W   R12,R10
						   56309 => x"6C",
						   56310 => x"92",		-- 00dbf6: 9212             CALL    &_lock
						   56311 => x"32",
						   56312 => x"F2",		-- 00dbf8: F220            
						   56313 => x"20",
						   56314 => x"0C",		-- 00dbfa: 0C4A             MOV.W   R10,R12
						   56315 => x"6A",
						   56316 => x"B0",		-- 00dbfc: B012             CALL    #strlen
						   56317 => x"32",
						   56318 => x"7A",		-- 00dbfe: 7AE1            
						   56319 => x"E1",
						   56320 => x"1F",		-- 00dc00: 1F43             MOV.W   #1,R15
						   56321 => x"63",
						   56322 => x"0F",		-- 00dc02: 0F5C             ADD.W   R12,R15
						   56323 => x"7C",
						   56324 => x"7C",		-- 00dc04: 7C40             MOV.B   #0x00f5,R12
						   56325 => x"60",
						   56326 => x"F5",		-- 00dc06: F500            
						   56327 => x"00",
						   56328 => x"3D",		-- 00dc08: 3D40             MOV.W   #0x219e,R13
						   56329 => x"60",
						   56330 => x"9E",		-- 00dc0a: 9E21            
						   56331 => x"21",
						   56332 => x"0E",		-- 00dc0c: 0E4A             MOV.W   R10,R14
						   56333 => x"6A",
						   56334 => x"B0",		-- 00dc0e: B012             CALL    #__TI_writemsg
						   56335 => x"32",
						   56336 => x"92",		-- 00dc10: 92DD            
						   56337 => x"DD",
						   56338 => x"3C",		-- 00dc12: 3C40             MOV.W   #0x219e,R12
						   56339 => x"60",
						   56340 => x"9E",		-- 00dc14: 9E21            
						   56341 => x"21",
						   56342 => x"0D",		-- 00dc16: 0D43             CLR.W   R13
						   56343 => x"63",
						   56344 => x"B0",		-- 00dc18: B012             CALL    #__TI_readmsg
						   56345 => x"32",
						   56346 => x"1C",		-- 00dc1a: 1CDE            
						   56347 => x"DE",
						   56348 => x"5F",		-- 00dc1c: 5F42             MOV.B   &parmbuf,R15
						   56349 => x"62",
						   56350 => x"9E",		-- 00dc1e: 9E21            
						   56351 => x"21",
						   56352 => x"5A",		-- 00dc20: 5A42             MOV.B   &0x219f,R10
						   56353 => x"62",
						   56354 => x"9F",		-- 00dc22: 9F21            
						   56355 => x"21",
						   56356 => x"8A",		-- 00dc24: 8A10             SWPB    R10
						   56357 => x"30",
						   56358 => x"0A",		-- 00dc26: 0A5F             ADD.W   R15,R10
						   56359 => x"7F",
						   56360 => x"92",		-- 00dc28: 9212             CALL    &_unlock
						   56361 => x"32",
						   56362 => x"F4",		-- 00dc2a: F420            
						   56363 => x"20",
						   56364 => x"0C",		-- 00dc2c: 0C4A             MOV.W   R10,R12
						   56365 => x"6A",
						   56366 => x"3A",		-- 00dc2e: 3A41             POP.W   R10
						   56367 => x"61",
						   56368 => x"30",		-- 00dc30: 3041             RET     
						   56369 => x"61",
						   -- Begin: __mspabi_divli
						   -- Begin: __mspabi_remli
						   56370 => x"0A",		-- 00dc32: 0A12             PUSH    R10
						   56371 => x"32",
						   56372 => x"0A",		-- 00dc34: 0A43             CLR.W   R10
						   56373 => x"63",
						   56374 => x"0F",		-- 00dc36: 0F93             TST.W   R15
						   56375 => x"B3",
						   56376 => x"05",		-- 00dc38: 0534             JGE     (dvd_sign)
						   56377 => x"54",
						   56378 => x"3E",		-- 00dc3a: 3EE3             INV.W   R14
						   56379 => x"03",
						   56380 => x"3F",		-- 00dc3c: 3FE3             INV.W   R15
						   56381 => x"03",
						   56382 => x"1E",		-- 00dc3e: 1E53             INC.W   R14
						   56383 => x"73",
						   56384 => x"0F",		-- 00dc40: 0F63             ADC.W   R15
						   56385 => x"83",
						   56386 => x"1A",		-- 00dc42: 1AD3             BIS.W   #1,R10
						   56387 => x"F3",
						   -- Begin: dvd_sign
						   56388 => x"0D",		-- 00dc44: 0D93             TST.W   R13
						   56389 => x"B3",
						   56390 => x"05",		-- 00dc46: 0534             JGE     (perform_divide)
						   56391 => x"54",
						   56392 => x"3C",		-- 00dc48: 3CE3             INV.W   R12
						   56393 => x"03",
						   56394 => x"3D",		-- 00dc4a: 3DE3             INV.W   R13
						   56395 => x"03",
						   56396 => x"1C",		-- 00dc4c: 1C53             INC.W   R12
						   56397 => x"73",
						   56398 => x"0D",		-- 00dc4e: 0D63             ADC.W   R13
						   56399 => x"83",
						   56400 => x"3A",		-- 00dc50: 3AE3             INV.W   R10
						   56401 => x"03",
						   -- Begin: perform_divide
						   56402 => x"B0",		-- 00dc52: B012             CALL    #__mspabi_divul
						   56403 => x"32",
						   56404 => x"7C",		-- 00dc54: 7CD8            
						   56405 => x"D8",
						   56406 => x"1A",		-- 00dc56: 1AB3             BIT.W   #1,R10
						   56407 => x"D3",
						   56408 => x"04",		-- 00dc58: 0424             JEQ     (rem_sign)
						   56409 => x"44",
						   56410 => x"3C",		-- 00dc5a: 3CE3             INV.W   R12
						   56411 => x"03",
						   56412 => x"3D",		-- 00dc5c: 3DE3             INV.W   R13
						   56413 => x"03",
						   56414 => x"1C",		-- 00dc5e: 1C53             INC.W   R12
						   56415 => x"73",
						   56416 => x"0D",		-- 00dc60: 0D63             ADC.W   R13
						   56417 => x"83",
						   -- Begin: rem_sign
						   56418 => x"2A",		-- 00dc62: 2AB3             BIT.W   #2,R10
						   56419 => x"D3",
						   56420 => x"04",		-- 00dc64: 0424             JEQ     (div_exit)
						   56421 => x"44",
						   56422 => x"3E",		-- 00dc66: 3EE3             INV.W   R14
						   56423 => x"03",
						   56424 => x"3F",		-- 00dc68: 3FE3             INV.W   R15
						   56425 => x"03",
						   56426 => x"1E",		-- 00dc6a: 1E53             INC.W   R14
						   56427 => x"73",
						   56428 => x"0F",		-- 00dc6c: 0F63             ADC.W   R15
						   56429 => x"83",
						   -- Begin: div_exit
						   56430 => x"3A",		-- 00dc6e: 3A41             POP.W   R10
						   56431 => x"61",
						   56432 => x"30",		-- 00dc70: 3041             RET     
						   56433 => x"61",
						   -- Begin: __mspabi_sral_15
						   56434 => x"0D",		-- 00dc72: 0D11             RRA     R13
						   56435 => x"31",
						   56436 => x"0C",		-- 00dc74: 0C10             RRC     R12
						   56437 => x"30",
						   -- Begin: __mspabi_sral_14
						   56438 => x"0D",		-- 00dc76: 0D11             RRA     R13
						   56439 => x"31",
						   56440 => x"0C",		-- 00dc78: 0C10             RRC     R12
						   56441 => x"30",
						   -- Begin: __mspabi_sral_13
						   56442 => x"0D",		-- 00dc7a: 0D11             RRA     R13
						   56443 => x"31",
						   56444 => x"0C",		-- 00dc7c: 0C10             RRC     R12
						   56445 => x"30",
						   -- Begin: __mspabi_sral_12
						   56446 => x"0D",		-- 00dc7e: 0D11             RRA     R13
						   56447 => x"31",
						   56448 => x"0C",		-- 00dc80: 0C10             RRC     R12
						   56449 => x"30",
						   -- Begin: __mspabi_sral_11
						   56450 => x"0D",		-- 00dc82: 0D11             RRA     R13
						   56451 => x"31",
						   56452 => x"0C",		-- 00dc84: 0C10             RRC     R12
						   56453 => x"30",
						   -- Begin: __mspabi_sral_10
						   56454 => x"0D",		-- 00dc86: 0D11             RRA     R13
						   56455 => x"31",
						   56456 => x"0C",		-- 00dc88: 0C10             RRC     R12
						   56457 => x"30",
						   -- Begin: __mspabi_sral_9
						   56458 => x"0D",		-- 00dc8a: 0D11             RRA     R13
						   56459 => x"31",
						   56460 => x"0C",		-- 00dc8c: 0C10             RRC     R12
						   56461 => x"30",
						   -- Begin: __mspabi_sral_8
						   56462 => x"0D",		-- 00dc8e: 0D11             RRA     R13
						   56463 => x"31",
						   56464 => x"0C",		-- 00dc90: 0C10             RRC     R12
						   56465 => x"30",
						   -- Begin: __mspabi_sral_7
						   56466 => x"0D",		-- 00dc92: 0D11             RRA     R13
						   56467 => x"31",
						   56468 => x"0C",		-- 00dc94: 0C10             RRC     R12
						   56469 => x"30",
						   -- Begin: __mspabi_sral_6
						   56470 => x"0D",		-- 00dc96: 0D11             RRA     R13
						   56471 => x"31",
						   56472 => x"0C",		-- 00dc98: 0C10             RRC     R12
						   56473 => x"30",
						   -- Begin: __mspabi_sral_5
						   56474 => x"0D",		-- 00dc9a: 0D11             RRA     R13
						   56475 => x"31",
						   56476 => x"0C",		-- 00dc9c: 0C10             RRC     R12
						   56477 => x"30",
						   -- Begin: __mspabi_sral_4
						   56478 => x"0D",		-- 00dc9e: 0D11             RRA     R13
						   56479 => x"31",
						   56480 => x"0C",		-- 00dca0: 0C10             RRC     R12
						   56481 => x"30",
						   -- Begin: __mspabi_sral_3
						   56482 => x"0D",		-- 00dca2: 0D11             RRA     R13
						   56483 => x"31",
						   56484 => x"0C",		-- 00dca4: 0C10             RRC     R12
						   56485 => x"30",
						   -- Begin: __mspabi_sral_2
						   56486 => x"0D",		-- 00dca6: 0D11             RRA     R13
						   56487 => x"31",
						   56488 => x"0C",		-- 00dca8: 0C10             RRC     R12
						   56489 => x"30",
						   -- Begin: __mspabi_sral_1
						   56490 => x"0D",		-- 00dcaa: 0D11             RRA     R13
						   56491 => x"31",
						   56492 => x"0C",		-- 00dcac: 0C10             RRC     R12
						   56493 => x"30",
						   56494 => x"30",		-- 00dcae: 3041             RET     
						   56495 => x"61",
						   -- Begin: __mspabi_slll_15
						   56496 => x"0C",		-- 00dcb0: 0C5C             RLA.W   R12
						   56497 => x"7C",
						   56498 => x"0D",		-- 00dcb2: 0D6D             RLC.W   R13
						   56499 => x"8D",
						   -- Begin: __mspabi_slll_14
						   56500 => x"0C",		-- 00dcb4: 0C5C             RLA.W   R12
						   56501 => x"7C",
						   56502 => x"0D",		-- 00dcb6: 0D6D             RLC.W   R13
						   56503 => x"8D",
						   -- Begin: __mspabi_slll_13
						   56504 => x"0C",		-- 00dcb8: 0C5C             RLA.W   R12
						   56505 => x"7C",
						   56506 => x"0D",		-- 00dcba: 0D6D             RLC.W   R13
						   56507 => x"8D",
						   -- Begin: __mspabi_slll_12
						   56508 => x"0C",		-- 00dcbc: 0C5C             RLA.W   R12
						   56509 => x"7C",
						   56510 => x"0D",		-- 00dcbe: 0D6D             RLC.W   R13
						   56511 => x"8D",
						   -- Begin: __mspabi_slll_11
						   56512 => x"0C",		-- 00dcc0: 0C5C             RLA.W   R12
						   56513 => x"7C",
						   56514 => x"0D",		-- 00dcc2: 0D6D             RLC.W   R13
						   56515 => x"8D",
						   -- Begin: __mspabi_slll_10
						   56516 => x"0C",		-- 00dcc4: 0C5C             RLA.W   R12
						   56517 => x"7C",
						   56518 => x"0D",		-- 00dcc6: 0D6D             RLC.W   R13
						   56519 => x"8D",
						   -- Begin: __mspabi_slll_9
						   56520 => x"0C",		-- 00dcc8: 0C5C             RLA.W   R12
						   56521 => x"7C",
						   56522 => x"0D",		-- 00dcca: 0D6D             RLC.W   R13
						   56523 => x"8D",
						   -- Begin: __mspabi_slll_8
						   56524 => x"0C",		-- 00dccc: 0C5C             RLA.W   R12
						   56525 => x"7C",
						   56526 => x"0D",		-- 00dcce: 0D6D             RLC.W   R13
						   56527 => x"8D",
						   -- Begin: __mspabi_slll_7
						   56528 => x"0C",		-- 00dcd0: 0C5C             RLA.W   R12
						   56529 => x"7C",
						   56530 => x"0D",		-- 00dcd2: 0D6D             RLC.W   R13
						   56531 => x"8D",
						   -- Begin: __mspabi_slll_6
						   56532 => x"0C",		-- 00dcd4: 0C5C             RLA.W   R12
						   56533 => x"7C",
						   56534 => x"0D",		-- 00dcd6: 0D6D             RLC.W   R13
						   56535 => x"8D",
						   -- Begin: __mspabi_slll_5
						   56536 => x"0C",		-- 00dcd8: 0C5C             RLA.W   R12
						   56537 => x"7C",
						   56538 => x"0D",		-- 00dcda: 0D6D             RLC.W   R13
						   56539 => x"8D",
						   -- Begin: __mspabi_slll_4
						   56540 => x"0C",		-- 00dcdc: 0C5C             RLA.W   R12
						   56541 => x"7C",
						   56542 => x"0D",		-- 00dcde: 0D6D             RLC.W   R13
						   56543 => x"8D",
						   -- Begin: __mspabi_slll_3
						   56544 => x"0C",		-- 00dce0: 0C5C             RLA.W   R12
						   56545 => x"7C",
						   56546 => x"0D",		-- 00dce2: 0D6D             RLC.W   R13
						   56547 => x"8D",
						   -- Begin: __mspabi_slll_2
						   56548 => x"0C",		-- 00dce4: 0C5C             RLA.W   R12
						   56549 => x"7C",
						   56550 => x"0D",		-- 00dce6: 0D6D             RLC.W   R13
						   56551 => x"8D",
						   -- Begin: __mspabi_slll_1
						   56552 => x"0C",		-- 00dce8: 0C5C             RLA.W   R12
						   56553 => x"7C",
						   56554 => x"0D",		-- 00dcea: 0D6D             RLC.W   R13
						   56555 => x"8D",
						   56556 => x"30",		-- 00dcec: 3041             RET     
						   56557 => x"61",
						   -- Begin: printf
						   56558 => x"0A",		-- 00dcee: 0A12             PUSH    R10
						   56559 => x"32",
						   56560 => x"21",		-- 00dcf0: 2183             DECD.W  SP
						   56561 => x"A3",
						   56562 => x"92",		-- 00dcf2: 9212             CALL    &_lock
						   56563 => x"32",
						   56564 => x"F2",		-- 00dcf4: F220            
						   56565 => x"20",
						   56566 => x"B2",		-- 00dcf6: B293             CMP.W   #-1,&0x200c
						   56567 => x"B3",
						   56568 => x"0C",		-- 00dcf8: 0C20            
						   56569 => x"20",
						   56570 => x"02",		-- 00dcfa: 0220             JNE     ($C$L1)
						   56571 => x"40",
						   56572 => x"3A",		-- 00dcfc: 3A43             MOV.W   #-1,R10
						   56573 => x"63",
						   56574 => x"0F",		-- 00dcfe: 0F3C             JMP     ($C$L2)
						   56575 => x"5C",
						   56576 => x"B1",		-- 00dd00: B140             MOV.W   #0xe1be,0x0000(SP)
						   56577 => x"60",
						   56578 => x"BE",		-- 00dd02: BEE1            
						   56579 => x"E1",
						   56580 => x"00",		-- 00dd04: 0000            
						   56581 => x"00",
						   56582 => x"0D",		-- 00dd06: 0D41             MOV.W   SP,R13
						   56583 => x"61",
						   56584 => x"3D",		-- 00dd08: 3D52             ADD.W   #8,R13
						   56585 => x"72",
						   56586 => x"3E",		-- 00dd0a: 3E40             MOV.W   #0x200c,R14
						   56587 => x"60",
						   56588 => x"0C",		-- 00dd0c: 0C20            
						   56589 => x"20",
						   56590 => x"0C",		-- 00dd0e: 0C41             MOV.W   SP,R12
						   56591 => x"61",
						   56592 => x"3C",		-- 00dd10: 3C50             ADD.W   #0x0006,R12
						   56593 => x"70",
						   56594 => x"06",		-- 00dd12: 0600            
						   56595 => x"00",
						   56596 => x"3F",		-- 00dd14: 3F40             MOV.W   #0xe1b2,R15
						   56597 => x"60",
						   56598 => x"B2",		-- 00dd16: B2E1            
						   56599 => x"E1",
						   56600 => x"B0",		-- 00dd18: B012             CALL    #__TI_printfi
						   56601 => x"32",
						   56602 => x"14",		-- 00dd1a: 14AC            
						   56603 => x"AC",
						   56604 => x"0A",		-- 00dd1c: 0A4C             MOV.W   R12,R10
						   56605 => x"6C",
						   56606 => x"92",		-- 00dd1e: 9212             CALL    &_unlock
						   56607 => x"32",
						   56608 => x"F4",		-- 00dd20: F420            
						   56609 => x"20",
						   56610 => x"0C",		-- 00dd22: 0C4A             MOV.W   R10,R12
						   56611 => x"6A",
						   56612 => x"21",		-- 00dd24: 2153             INCD.W  SP
						   56613 => x"73",
						   56614 => x"3A",		-- 00dd26: 3A41             POP.W   R10
						   56615 => x"61",
						   56616 => x"30",		-- 00dd28: 3041             RET     
						   56617 => x"61",
						   -- Begin: __TI_cleanup
						   56618 => x"0A",		-- 00dd2a: 0A12             PUSH    R10
						   56619 => x"32",
						   56620 => x"09",		-- 00dd2c: 0912             PUSH    R9
						   56621 => x"32",
						   56622 => x"3C",		-- 00dd2e: 3C40             MOV.W   #0x2000,R12
						   56623 => x"60",
						   56624 => x"00",		-- 00dd30: 0020            
						   56625 => x"20",
						   56626 => x"B0",		-- 00dd32: B012             CALL    #__TI_closefile
						   56627 => x"32",
						   56628 => x"18",		-- 00dd34: 18D4            
						   56629 => x"D4",
						   56630 => x"A2",		-- 00dd36: A293             CMP.W   #2,&__TI_ft_end
						   56631 => x"B3",
						   56632 => x"F6",		-- 00dd38: F620            
						   56633 => x"20",
						   56634 => x"0F",		-- 00dd3a: 0F38             JL      ($C$L37)
						   56635 => x"58",
						   56636 => x"3A",		-- 00dd3c: 3A40             MOV.W   #0x200c,R10
						   56637 => x"60",
						   56638 => x"0C",		-- 00dd3e: 0C20            
						   56639 => x"20",
						   56640 => x"19",		-- 00dd40: 1943             MOV.W   #1,R9
						   56641 => x"63",
						   56642 => x"8A",		-- 00dd42: 8A93             TST.W   0x0000(R10)
						   56643 => x"B3",
						   56644 => x"00",		-- 00dd44: 0000            
						   56645 => x"00",
						   56646 => x"03",		-- 00dd46: 0338             JL      ($C$L36)
						   56647 => x"58",
						   56648 => x"0C",		-- 00dd48: 0C4A             MOV.W   R10,R12
						   56649 => x"6A",
						   56650 => x"B0",		-- 00dd4a: B012             CALL    #__TI_closefile
						   56651 => x"32",
						   56652 => x"18",		-- 00dd4c: 18D4            
						   56653 => x"D4",
						   56654 => x"3A",		-- 00dd4e: 3A50             ADD.W   #0x000c,R10
						   56655 => x"70",
						   56656 => x"0C",		-- 00dd50: 0C00            
						   56657 => x"00",
						   56658 => x"19",		-- 00dd52: 1953             INC.W   R9
						   56659 => x"73",
						   56660 => x"19",		-- 00dd54: 1992             CMP.W   &__TI_ft_end,R9
						   56661 => x"B2",
						   56662 => x"F6",		-- 00dd56: F620            
						   56663 => x"20",
						   56664 => x"F4",		-- 00dd58: F43B             JL      ($C$L35)
						   56665 => x"5B",
						   56666 => x"30",		-- 00dd5a: 3040             BR      #__mspabi_func_epilog_2
						   56667 => x"60",
						   56668 => x"64",		-- 00dd5c: 64E1            
						   56669 => x"E1",
						   -- Begin: finddevice
						   56670 => x"0A",		-- 00dd5e: 0A12             PUSH    R10
						   56671 => x"32",
						   56672 => x"09",		-- 00dd60: 0912             PUSH    R9
						   56673 => x"32",
						   56674 => x"08",		-- 00dd62: 0812             PUSH    R8
						   56675 => x"32",
						   56676 => x"08",		-- 00dd64: 084C             MOV.W   R12,R8
						   56677 => x"6C",
						   56678 => x"C8",		-- 00dd66: C893             TST.B   0x0000(R8)
						   56679 => x"B3",
						   56680 => x"00",		-- 00dd68: 0000            
						   56681 => x"00",
						   56682 => x"10",		-- 00dd6a: 1024             JEQ     ($C$L3)
						   56683 => x"44",
						   56684 => x"3A",		-- 00dd6c: 3A40             MOV.W   #0x2092,R10
						   56685 => x"60",
						   56686 => x"92",		-- 00dd6e: 9220            
						   56687 => x"20",
						   56688 => x"29",		-- 00dd70: 2943             MOV.W   #2,R9
						   56689 => x"63",
						   56690 => x"0C",		-- 00dd72: 0C4A             MOV.W   R10,R12
						   56691 => x"6A",
						   56692 => x"0D",		-- 00dd74: 0D48             MOV.W   R8,R13
						   56693 => x"68",
						   56694 => x"B0",		-- 00dd76: B012             CALL    #strcmp
						   56695 => x"32",
						   56696 => x"92",		-- 00dd78: 92E0            
						   56697 => x"E0",
						   56698 => x"0C",		-- 00dd7a: 0C93             TST.W   R12
						   56699 => x"B3",
						   56700 => x"03",		-- 00dd7c: 0320             JNE     ($C$L2)
						   56701 => x"40",
						   56702 => x"0C",		-- 00dd7e: 0C4A             MOV.W   R10,R12
						   56703 => x"6A",
						   56704 => x"30",		-- 00dd80: 3040             BR      #__mspabi_func_epilog_3
						   56705 => x"60",
						   56706 => x"62",		-- 00dd82: 62E1            
						   56707 => x"E1",
						   56708 => x"3A",		-- 00dd84: 3A50             ADD.W   #0x001a,R10
						   56709 => x"70",
						   56710 => x"1A",		-- 00dd86: 1A00            
						   56711 => x"00",
						   56712 => x"19",		-- 00dd88: 1983             DEC.W   R9
						   56713 => x"A3",
						   56714 => x"F3",		-- 00dd8a: F323             JNE     ($C$L1)
						   56715 => x"43",
						   56716 => x"0C",		-- 00dd8c: 0C43             CLR.W   R12
						   56717 => x"63",
						   56718 => x"30",		-- 00dd8e: 3040             BR      #__mspabi_func_epilog_3
						   56719 => x"60",
						   56720 => x"62",		-- 00dd90: 62E1            
						   56721 => x"E1",
						   -- Begin: __TI_writemsg
						   56722 => x"82",		-- 00dd92: 824F             MOV.W   R15,&_CIOBUF_
						   56723 => x"6F",
						   56724 => x"00",		-- 00dd94: 0080            
						   56725 => x"80",
						   56726 => x"C2",		-- 00dd96: C24C             MOV.B   R12,&0x8002
						   56727 => x"6C",
						   56728 => x"02",		-- 00dd98: 0280            
						   56729 => x"80",
						   56730 => x"3C",		-- 00dd9a: 3C40             MOV.W   #0x8003,R12
						   56731 => x"60",
						   56732 => x"03",		-- 00dd9c: 0380            
						   56733 => x"80",
						   56734 => x"3B",		-- 00dd9e: 3B42             MOV.W   #8,R11
						   56735 => x"62",
						   56736 => x"1C",		-- 00dda0: 1C53             INC.W   R12
						   56737 => x"73",
						   56738 => x"FC",		-- 00dda2: FC4D             MOV.B   @R13+,0xffff(R12)
						   56739 => x"6D",
						   56740 => x"FF",		-- 00dda4: FFFF            
						   56741 => x"FF",
						   56742 => x"1B",		-- 00dda6: 1B83             DEC.W   R11
						   56743 => x"A3",
						   56744 => x"FB",		-- 00dda8: FB23             JNE     ($C$L1)
						   56745 => x"43",
						   56746 => x"0F",		-- 00ddaa: 0F93             TST.W   R15
						   56747 => x"B3",
						   56748 => x"07",		-- 00ddac: 0724             JEQ     (C$$IO$$)
						   56749 => x"44",
						   56750 => x"3D",		-- 00ddae: 3D40             MOV.W   #0x800b,R13
						   56751 => x"60",
						   56752 => x"0B",		-- 00ddb0: 0B80            
						   56753 => x"80",
						   56754 => x"1D",		-- 00ddb2: 1D53             INC.W   R13
						   56755 => x"73",
						   56756 => x"FD",		-- 00ddb4: FD4E             MOV.B   @R14+,0xffff(R13)
						   56757 => x"6E",
						   56758 => x"FF",		-- 00ddb6: FFFF            
						   56759 => x"FF",
						   56760 => x"1F",		-- 00ddb8: 1F83             DEC.W   R15
						   56761 => x"A3",
						   56762 => x"FB",		-- 00ddba: FB23             JNE     ($C$L2)
						   56763 => x"43",
						   56764 => x"03",		-- 00ddbc: 0343             NOP     
						   56765 => x"63",
						   56766 => x"30",		-- 00ddbe: 3041             RET     
						   56767 => x"61",
						   -- Begin: __mspabi_subd
						   56768 => x"31",		-- 00ddc0: 3182             SUB.W   #8,SP
						   56769 => x"A2",
						   56770 => x"81",		-- 00ddc2: 814C             MOV.W   R12,0x0000(SP)
						   56771 => x"6C",
						   56772 => x"00",		-- 00ddc4: 0000            
						   56773 => x"00",
						   56774 => x"81",		-- 00ddc6: 814D             MOV.W   R13,0x0002(SP)
						   56775 => x"6D",
						   56776 => x"02",		-- 00ddc8: 0200            
						   56777 => x"00",
						   56778 => x"81",		-- 00ddca: 814E             MOV.W   R14,0x0004(SP)
						   56779 => x"6E",
						   56780 => x"04",		-- 00ddcc: 0400            
						   56781 => x"00",
						   56782 => x"81",		-- 00ddce: 814F             MOV.W   R15,0x0006(SP)
						   56783 => x"6F",
						   56784 => x"06",		-- 00ddd0: 0600            
						   56785 => x"00",
						   56786 => x"F1",		-- 00ddd2: F1E0             XOR.B   #0x0080,0x0007(SP)
						   56787 => x"00",
						   56788 => x"80",		-- 00ddd4: 8000            
						   56789 => x"00",
						   56790 => x"07",		-- 00ddd6: 0700            
						   56791 => x"00",
						   56792 => x"2C",		-- 00ddd8: 2C41             MOV.W   @SP,R12
						   56793 => x"61",
						   56794 => x"1D",		-- 00ddda: 1D41             MOV.W   0x0002(SP),R13
						   56795 => x"61",
						   56796 => x"02",		-- 00dddc: 0200            
						   56797 => x"00",
						   56798 => x"1E",		-- 00ddde: 1E41             MOV.W   0x0004(SP),R14
						   56799 => x"61",
						   56800 => x"04",		-- 00dde0: 0400            
						   56801 => x"00",
						   56802 => x"1F",		-- 00dde2: 1F41             MOV.W   0x0006(SP),R15
						   56803 => x"61",
						   56804 => x"06",		-- 00dde4: 0600            
						   56805 => x"00",
						   56806 => x"B0",		-- 00dde6: B012             CALL    #__mspabi_addd
						   56807 => x"32",
						   56808 => x"46",		-- 00dde8: 469A            
						   56809 => x"9A",
						   56810 => x"31",		-- 00ddea: 3152             ADD.W   #8,SP
						   56811 => x"72",
						   56812 => x"30",		-- 00ddec: 3041             RET     
						   56813 => x"61",
						   -- Begin: copysignl
						   -- Begin: copysign
						   56814 => x"0A",		-- 00ddee: 0A12             PUSH    R10
						   56815 => x"32",
						   56816 => x"1A",		-- 00ddf0: 1A41             MOV.W   0x0008(SP),R10
						   56817 => x"61",
						   56818 => x"08",		-- 00ddf2: 0800            
						   56819 => x"00",
						   56820 => x"1B",		-- 00ddf4: 1B41             MOV.W   0x000a(SP),R11
						   56821 => x"61",
						   56822 => x"0A",		-- 00ddf6: 0A00            
						   56823 => x"00",
						   56824 => x"0A",		-- 00ddf8: 0AF3             AND.W   #0,R10
						   56825 => x"13",
						   56826 => x"3B",		-- 00ddfa: 3BF0             AND.W   #0x8000,R11
						   56827 => x"10",
						   56828 => x"00",		-- 00ddfc: 0080            
						   56829 => x"80",
						   56830 => x"3E",		-- 00ddfe: 3EF3             AND.W   #-1,R14
						   56831 => x"13",
						   56832 => x"3F",		-- 00de00: 3FF0             AND.W   #0x7fff,R15
						   56833 => x"10",
						   56834 => x"FF",		-- 00de02: FF7F            
						   56835 => x"7F",
						   56836 => x"0E",		-- 00de04: 0EDA             BIS.W   R10,R14
						   56837 => x"FA",
						   56838 => x"0F",		-- 00de06: 0FDB             BIS.W   R11,R15
						   56839 => x"FB",
						   56840 => x"0B",		-- 00de08: 0B43             CLR.W   R11
						   56841 => x"63",
						   56842 => x"0B",		-- 00de0a: 0BDD             BIS.W   R13,R11
						   56843 => x"FD",
						   56844 => x"0D",		-- 00de0c: 0D43             CLR.W   R13
						   56845 => x"63",
						   56846 => x"0D",		-- 00de0e: 0DDC             BIS.W   R12,R13
						   56847 => x"FC",
						   56848 => x"0E",		-- 00de10: 0ED3             BIS.W   #0,R14
						   56849 => x"F3",
						   56850 => x"0F",		-- 00de12: 0FD3             BIS.W   #0,R15
						   56851 => x"F3",
						   56852 => x"0C",		-- 00de14: 0C4D             MOV.W   R13,R12
						   56853 => x"6D",
						   56854 => x"0D",		-- 00de16: 0D4B             MOV.W   R11,R13
						   56855 => x"6B",
						   56856 => x"3A",		-- 00de18: 3A41             POP.W   R10
						   56857 => x"61",
						   56858 => x"30",		-- 00de1a: 3041             RET     
						   56859 => x"61",
						   -- Begin: __TI_readmsg
						   56860 => x"1F",		-- 00de1c: 1F42             MOV.W   &_CIOBUF_,R15
						   56861 => x"62",
						   56862 => x"00",		-- 00de1e: 0080            
						   56863 => x"80",
						   56864 => x"3B",		-- 00de20: 3B40             MOV.W   #0x8002,R11
						   56865 => x"60",
						   56866 => x"02",		-- 00de22: 0280            
						   56867 => x"80",
						   56868 => x"3E",		-- 00de24: 3E42             MOV.W   #8,R14
						   56869 => x"62",
						   56870 => x"1C",		-- 00de26: 1C53             INC.W   R12
						   56871 => x"73",
						   56872 => x"FC",		-- 00de28: FC4B             MOV.B   @R11+,0xffff(R12)
						   56873 => x"6B",
						   56874 => x"FF",		-- 00de2a: FFFF            
						   56875 => x"FF",
						   56876 => x"1E",		-- 00de2c: 1E83             DEC.W   R14
						   56877 => x"A3",
						   56878 => x"FB",		-- 00de2e: FB23             JNE     ($C$L4)
						   56879 => x"43",
						   56880 => x"0D",		-- 00de30: 0D93             TST.W   R13
						   56881 => x"B3",
						   56882 => x"09",		-- 00de32: 0924             JEQ     ($C$L6)
						   56883 => x"44",
						   56884 => x"0F",		-- 00de34: 0F93             TST.W   R15
						   56885 => x"B3",
						   56886 => x"07",		-- 00de36: 0724             JEQ     ($C$L6)
						   56887 => x"44",
						   56888 => x"3E",		-- 00de38: 3E40             MOV.W   #0x800a,R14
						   56889 => x"60",
						   56890 => x"0A",		-- 00de3a: 0A80            
						   56891 => x"80",
						   56892 => x"1D",		-- 00de3c: 1D53             INC.W   R13
						   56893 => x"73",
						   56894 => x"FD",		-- 00de3e: FD4E             MOV.B   @R14+,0xffff(R13)
						   56895 => x"6E",
						   56896 => x"FF",		-- 00de40: FFFF            
						   56897 => x"FF",
						   56898 => x"1F",		-- 00de42: 1F83             DEC.W   R15
						   56899 => x"A3",
						   56900 => x"FB",		-- 00de44: FB23             JNE     ($C$L5)
						   56901 => x"43",
						   56902 => x"30",		-- 00de46: 3041             RET     
						   56903 => x"61",
						   -- Begin: __mspabi_srai
						   56904 => x"3D",		-- 00de48: 3DF0             AND.W   #0x000f,R13
						   56905 => x"10",
						   56906 => x"0F",		-- 00de4a: 0F00            
						   56907 => x"00",
						   56908 => x"3D",		-- 00de4c: 3DE0             XOR.W   #0x000f,R13
						   56909 => x"00",
						   56910 => x"0F",		-- 00de4e: 0F00            
						   56911 => x"00",
						   56912 => x"0D",		-- 00de50: 0D5D             RLA.W   R13
						   56913 => x"7D",
						   56914 => x"00",		-- 00de52: 005D             ADD.W   R13,PC
						   56915 => x"7D",
						   -- Begin: __mspabi_srai_15
						   56916 => x"0C",		-- 00de54: 0C11             RRA     R12
						   56917 => x"31",
						   -- Begin: __mspabi_srai_14
						   56918 => x"0C",		-- 00de56: 0C11             RRA     R12
						   56919 => x"31",
						   -- Begin: __mspabi_srai_13
						   56920 => x"0C",		-- 00de58: 0C11             RRA     R12
						   56921 => x"31",
						   -- Begin: __mspabi_srai_12
						   56922 => x"0C",		-- 00de5a: 0C11             RRA     R12
						   56923 => x"31",
						   -- Begin: __mspabi_srai_11
						   56924 => x"0C",		-- 00de5c: 0C11             RRA     R12
						   56925 => x"31",
						   -- Begin: __mspabi_srai_10
						   56926 => x"0C",		-- 00de5e: 0C11             RRA     R12
						   56927 => x"31",
						   -- Begin: __mspabi_srai_9
						   56928 => x"0C",		-- 00de60: 0C11             RRA     R12
						   56929 => x"31",
						   -- Begin: __mspabi_srai_8
						   56930 => x"0C",		-- 00de62: 0C11             RRA     R12
						   56931 => x"31",
						   -- Begin: __mspabi_srai_7
						   56932 => x"0C",		-- 00de64: 0C11             RRA     R12
						   56933 => x"31",
						   -- Begin: __mspabi_srai_6
						   56934 => x"0C",		-- 00de66: 0C11             RRA     R12
						   56935 => x"31",
						   -- Begin: __mspabi_srai_5
						   56936 => x"0C",		-- 00de68: 0C11             RRA     R12
						   56937 => x"31",
						   -- Begin: __mspabi_srai_4
						   56938 => x"0C",		-- 00de6a: 0C11             RRA     R12
						   56939 => x"31",
						   -- Begin: __mspabi_srai_3
						   56940 => x"0C",		-- 00de6c: 0C11             RRA     R12
						   56941 => x"31",
						   -- Begin: __mspabi_srai_2
						   56942 => x"0C",		-- 00de6e: 0C11             RRA     R12
						   56943 => x"31",
						   -- Begin: __mspabi_srai_1
						   56944 => x"0C",		-- 00de70: 0C11             RRA     R12
						   56945 => x"31",
						   56946 => x"30",		-- 00de72: 3041             RET     
						   56947 => x"61",
						   -- Begin: __mspabi_slli
						   56948 => x"3D",		-- 00de74: 3DF0             AND.W   #0x000f,R13
						   56949 => x"10",
						   56950 => x"0F",		-- 00de76: 0F00            
						   56951 => x"00",
						   56952 => x"3D",		-- 00de78: 3DE0             XOR.W   #0x000f,R13
						   56953 => x"00",
						   56954 => x"0F",		-- 00de7a: 0F00            
						   56955 => x"00",
						   56956 => x"0D",		-- 00de7c: 0D5D             RLA.W   R13
						   56957 => x"7D",
						   56958 => x"00",		-- 00de7e: 005D             ADD.W   R13,PC
						   56959 => x"7D",
						   -- Begin: __mspabi_slli_15
						   56960 => x"0C",		-- 00de80: 0C5C             RLA.W   R12
						   56961 => x"7C",
						   -- Begin: __mspabi_slli_14
						   56962 => x"0C",		-- 00de82: 0C5C             RLA.W   R12
						   56963 => x"7C",
						   -- Begin: __mspabi_slli_13
						   56964 => x"0C",		-- 00de84: 0C5C             RLA.W   R12
						   56965 => x"7C",
						   -- Begin: __mspabi_slli_12
						   56966 => x"0C",		-- 00de86: 0C5C             RLA.W   R12
						   56967 => x"7C",
						   -- Begin: __mspabi_slli_11
						   56968 => x"0C",		-- 00de88: 0C5C             RLA.W   R12
						   56969 => x"7C",
						   -- Begin: __mspabi_slli_10
						   56970 => x"0C",		-- 00de8a: 0C5C             RLA.W   R12
						   56971 => x"7C",
						   -- Begin: __mspabi_slli_9
						   56972 => x"0C",		-- 00de8c: 0C5C             RLA.W   R12
						   56973 => x"7C",
						   -- Begin: __mspabi_slli_8
						   56974 => x"0C",		-- 00de8e: 0C5C             RLA.W   R12
						   56975 => x"7C",
						   -- Begin: __mspabi_slli_7
						   56976 => x"0C",		-- 00de90: 0C5C             RLA.W   R12
						   56977 => x"7C",
						   -- Begin: __mspabi_slli_6
						   56978 => x"0C",		-- 00de92: 0C5C             RLA.W   R12
						   56979 => x"7C",
						   -- Begin: __mspabi_slli_5
						   56980 => x"0C",		-- 00de94: 0C5C             RLA.W   R12
						   56981 => x"7C",
						   -- Begin: __mspabi_slli_4
						   56982 => x"0C",		-- 00de96: 0C5C             RLA.W   R12
						   56983 => x"7C",
						   -- Begin: __mspabi_slli_3
						   56984 => x"0C",		-- 00de98: 0C5C             RLA.W   R12
						   56985 => x"7C",
						   -- Begin: __mspabi_slli_2
						   56986 => x"0C",		-- 00de9a: 0C5C             RLA.W   R12
						   56987 => x"7C",
						   -- Begin: __mspabi_slli_1
						   56988 => x"0C",		-- 00de9c: 0C5C             RLA.W   R12
						   56989 => x"7C",
						   56990 => x"30",		-- 00de9e: 3041             RET     
						   56991 => x"61",
						   -- Begin: strncpy
						   56992 => x"0E",		-- 00dea0: 0E93             TST.W   R14
						   56993 => x"B3",
						   56994 => x"13",		-- 00dea2: 1324             JEQ     ($C$L4)
						   56995 => x"44",
						   56996 => x"0F",		-- 00dea4: 0F4C             MOV.W   R12,R15
						   56997 => x"6C",
						   56998 => x"6B",		-- 00dea6: 6B4D             MOV.B   @R13,R11
						   56999 => x"6D",
						   57000 => x"1F",		-- 00dea8: 1F53             INC.W   R15
						   57001 => x"73",
						   57002 => x"CF",		-- 00deaa: CF4B             MOV.B   R11,0xffff(R15)
						   57003 => x"6B",
						   57004 => x"FF",		-- 00deac: FFFF            
						   57005 => x"FF",
						   57006 => x"0B",		-- 00deae: 0B93             TST.W   R11
						   57007 => x"B3",
						   57008 => x"03",		-- 00deb0: 0324             JEQ     ($C$L2)
						   57009 => x"44",
						   57010 => x"1D",		-- 00deb2: 1D53             INC.W   R13
						   57011 => x"73",
						   57012 => x"1E",		-- 00deb4: 1E83             DEC.W   R14
						   57013 => x"A3",
						   57014 => x"F7",		-- 00deb6: F723             JNE     ($C$L1)
						   57015 => x"43",
						   57016 => x"0D",		-- 00deb8: 0D4E             MOV.W   R14,R13
						   57017 => x"6E",
						   57018 => x"1E",		-- 00deba: 1E83             DEC.W   R14
						   57019 => x"A3",
						   57020 => x"2D",		-- 00debc: 2D93             CMP.W   #2,R13
						   57021 => x"B3",
						   57022 => x"05",		-- 00debe: 0528             JLO     ($C$L4)
						   57023 => x"48",
						   57024 => x"1F",		-- 00dec0: 1F53             INC.W   R15
						   57025 => x"73",
						   57026 => x"CF",		-- 00dec2: CF43             CLR.B   0xffff(R15)
						   57027 => x"63",
						   57028 => x"FF",		-- 00dec4: FFFF            
						   57029 => x"FF",
						   57030 => x"1E",		-- 00dec6: 1E83             DEC.W   R14
						   57031 => x"A3",
						   57032 => x"FB",		-- 00dec8: FB23             JNE     ($C$L3)
						   57033 => x"43",
						   57034 => x"30",		-- 00deca: 3041             RET     
						   57035 => x"61",
						   -- Begin: __mspabi_negd
						   57036 => x"31",		-- 00decc: 3182             SUB.W   #8,SP
						   57037 => x"A2",
						   57038 => x"81",		-- 00dece: 814C             MOV.W   R12,0x0000(SP)
						   57039 => x"6C",
						   57040 => x"00",		-- 00ded0: 0000            
						   57041 => x"00",
						   57042 => x"81",		-- 00ded2: 814D             MOV.W   R13,0x0002(SP)
						   57043 => x"6D",
						   57044 => x"02",		-- 00ded4: 0200            
						   57045 => x"00",
						   57046 => x"81",		-- 00ded6: 814E             MOV.W   R14,0x0004(SP)
						   57047 => x"6E",
						   57048 => x"04",		-- 00ded8: 0400            
						   57049 => x"00",
						   57050 => x"81",		-- 00deda: 814F             MOV.W   R15,0x0006(SP)
						   57051 => x"6F",
						   57052 => x"06",		-- 00dedc: 0600            
						   57053 => x"00",
						   57054 => x"F1",		-- 00dede: F1E0             XOR.B   #0x0080,0x0007(SP)
						   57055 => x"00",
						   57056 => x"80",		-- 00dee0: 8000            
						   57057 => x"00",
						   57058 => x"07",		-- 00dee2: 0700            
						   57059 => x"00",
						   57060 => x"2C",		-- 00dee4: 2C41             MOV.W   @SP,R12
						   57061 => x"61",
						   57062 => x"1D",		-- 00dee6: 1D41             MOV.W   0x0002(SP),R13
						   57063 => x"61",
						   57064 => x"02",		-- 00dee8: 0200            
						   57065 => x"00",
						   57066 => x"1E",		-- 00deea: 1E41             MOV.W   0x0004(SP),R14
						   57067 => x"61",
						   57068 => x"04",		-- 00deec: 0400            
						   57069 => x"00",
						   57070 => x"1F",		-- 00deee: 1F41             MOV.W   0x0006(SP),R15
						   57071 => x"61",
						   57072 => x"06",		-- 00def0: 0600            
						   57073 => x"00",
						   57074 => x"31",		-- 00def2: 3152             ADD.W   #8,SP
						   57075 => x"72",
						   57076 => x"30",		-- 00def4: 3041             RET     
						   57077 => x"61",
						   -- Begin: __mspabi_fixdi
						   57078 => x"B0",		-- 00def6: B012             CALL    #__mspabi_fixdli
						   57079 => x"32",
						   57080 => x"8A",		-- 00def8: 8AD4            
						   57081 => x"D4",
						   57082 => x"0D",		-- 00defa: 0D93             TST.W   R13
						   57083 => x"B3",
						   57084 => x"07",		-- 00defc: 0738             JL      ($C$L7)
						   57085 => x"58",
						   57086 => x"03",		-- 00defe: 0320             JNE     ($C$L6)
						   57087 => x"40",
						   57088 => x"3C",		-- 00df00: 3C90             CMP.W   #0x8000,R12
						   57089 => x"B0",
						   57090 => x"00",		-- 00df02: 0080            
						   57091 => x"80",
						   57092 => x"03",		-- 00df04: 0328             JLO     ($C$L7)
						   57093 => x"48",
						   57094 => x"3C",		-- 00df06: 3C40             MOV.W   #0x7fff,R12
						   57095 => x"60",
						   57096 => x"FF",		-- 00df08: FF7F            
						   57097 => x"7F",
						   57098 => x"30",		-- 00df0a: 3041             RET     
						   57099 => x"61",
						   57100 => x"3D",		-- 00df0c: 3D93             CMP.W   #-1,R13
						   57101 => x"B3",
						   57102 => x"04",		-- 00df0e: 0438             JL      ($C$L8)
						   57103 => x"58",
						   57104 => x"05",		-- 00df10: 0520             JNE     ($C$L9)
						   57105 => x"40",
						   57106 => x"3C",		-- 00df12: 3C90             CMP.W   #0x8000,R12
						   57107 => x"B0",
						   57108 => x"00",		-- 00df14: 0080            
						   57109 => x"80",
						   57110 => x"02",		-- 00df16: 022C             JHS     ($C$L9)
						   57111 => x"4C",
						   57112 => x"3C",		-- 00df18: 3C40             MOV.W   #0x8000,R12
						   57113 => x"60",
						   57114 => x"00",		-- 00df1a: 0080            
						   57115 => x"80",
						   57116 => x"30",		-- 00df1c: 3041             RET     
						   57117 => x"61",
						   -- Begin: free_list_insert
						   57118 => x"2F",		-- 00df1e: 2F4C             MOV.W   @R12,R15
						   57119 => x"6C",
						   57120 => x"1F",		-- 00df20: 1FC3             BIC.W   #1,R15
						   57121 => x"E3",
						   57122 => x"3E",		-- 00df22: 3E40             MOV.W   #0x21a6,R14
						   57123 => x"60",
						   57124 => x"A6",		-- 00df24: A621            
						   57125 => x"21",
						   57126 => x"03",		-- 00df26: 033C             JMP     ($C$L5)
						   57127 => x"5C",
						   57128 => x"2D",		-- 00df28: 2D42             MOV.W   #4,R13
						   57129 => x"62",
						   57130 => x"2D",		-- 00df2a: 2D5E             ADD.W   @R14,R13
						   57131 => x"7E",
						   57132 => x"0E",		-- 00df2c: 0E4D             MOV.W   R13,R14
						   57133 => x"6D",
						   57134 => x"2D",		-- 00df2e: 2D4E             MOV.W   @R14,R13
						   57135 => x"6E",
						   57136 => x"0D",		-- 00df30: 0D93             TST.W   R13
						   57137 => x"B3",
						   57138 => x"04",		-- 00df32: 0424             JEQ     ($C$L6)
						   57139 => x"44",
						   57140 => x"2D",		-- 00df34: 2D4D             MOV.W   @R13,R13
						   57141 => x"6D",
						   57142 => x"1D",		-- 00df36: 1DC3             BIC.W   #1,R13
						   57143 => x"E3",
						   57144 => x"0D",		-- 00df38: 0D9F             CMP.W   R15,R13
						   57145 => x"BF",
						   57146 => x"F6",		-- 00df3a: F62B             JLO     ($C$L4)
						   57147 => x"4B",
						   57148 => x"AC",		-- 00df3c: AC4E             MOV.W   @R14,0x0004(R12)
						   57149 => x"6E",
						   57150 => x"04",		-- 00df3e: 0400            
						   57151 => x"00",
						   57152 => x"8E",		-- 00df40: 8E4C             MOV.W   R12,0x0000(R14)
						   57153 => x"6C",
						   57154 => x"00",		-- 00df42: 0000            
						   57155 => x"00",
						   57156 => x"30",		-- 00df44: 3041             RET     
						   57157 => x"61",
						   -- Begin: remove
						   -- Begin: unlink
						   57158 => x"0A",		-- 00df46: 0A12             PUSH    R10
						   57159 => x"32",
						   57160 => x"21",		-- 00df48: 2183             DECD.W  SP
						   57161 => x"A3",
						   57162 => x"81",		-- 00df4a: 814C             MOV.W   R12,0x0000(SP)
						   57163 => x"6C",
						   57164 => x"00",		-- 00df4c: 0000            
						   57165 => x"00",
						   57166 => x"92",		-- 00df4e: 9212             CALL    &_lock
						   57167 => x"32",
						   57168 => x"F2",		-- 00df50: F220            
						   57169 => x"20",
						   57170 => x"0C",		-- 00df52: 0C41             MOV.W   SP,R12
						   57171 => x"61",
						   57172 => x"B0",		-- 00df54: B012             CALL    #getdevice
						   57173 => x"32",
						   57174 => x"24",		-- 00df56: 24D8            
						   57175 => x"D8",
						   57176 => x"0F",		-- 00df58: 0F4C             MOV.W   R12,R15
						   57177 => x"6C",
						   57178 => x"2C",		-- 00df5a: 2C41             MOV.W   @SP,R12
						   57179 => x"61",
						   57180 => x"9F",		-- 00df5c: 9F12             CALL    0x0016(R15)
						   57181 => x"32",
						   57182 => x"16",		-- 00df5e: 1600            
						   57183 => x"00",
						   57184 => x"0A",		-- 00df60: 0A4C             MOV.W   R12,R10
						   57185 => x"6C",
						   57186 => x"92",		-- 00df62: 9212             CALL    &_unlock
						   57187 => x"32",
						   57188 => x"F4",		-- 00df64: F420            
						   57189 => x"20",
						   57190 => x"0C",		-- 00df66: 0C4A             MOV.W   R10,R12
						   57191 => x"6A",
						   57192 => x"21",		-- 00df68: 2153             INCD.W  SP
						   57193 => x"73",
						   57194 => x"3A",		-- 00df6a: 3A41             POP.W   R10
						   57195 => x"61",
						   57196 => x"30",		-- 00df6c: 3041             RET     
						   57197 => x"61",
						   -- Begin: lseek
						   57198 => x"0C",		-- 00df6e: 0C93             TST.W   R12
						   57199 => x"B3",
						   57200 => x"0E",		-- 00df70: 0E38             JL      ($C$L1)
						   57201 => x"58",
						   57202 => x"3C",		-- 00df72: 3C90             CMP.W   #0x000a,R12
						   57203 => x"B0",
						   57204 => x"0A",		-- 00df74: 0A00            
						   57205 => x"00",
						   57206 => x"0B",		-- 00df76: 0B34             JGE     ($C$L1)
						   57207 => x"54",
						   57208 => x"0C",		-- 00df78: 0C5C             RLA.W   R12
						   57209 => x"7C",
						   57210 => x"0C",		-- 00df7a: 0C5C             RLA.W   R12
						   57211 => x"7C",
						   57212 => x"3C",		-- 00df7c: 3C50             ADD.W   #0x20c6,R12
						   57213 => x"70",
						   57214 => x"C6",		-- 00df7e: C620            
						   57215 => x"20",
						   57216 => x"2B",		-- 00df80: 2B4C             MOV.W   @R12,R11
						   57217 => x"6C",
						   57218 => x"0B",		-- 00df82: 0B93             TST.W   R11
						   57219 => x"B3",
						   57220 => x"04",		-- 00df84: 0424             JEQ     ($C$L1)
						   57221 => x"44",
						   57222 => x"1C",		-- 00df86: 1C4C             MOV.W   0x0002(R12),R12
						   57223 => x"6C",
						   57224 => x"02",		-- 00df88: 0200            
						   57225 => x"00",
						   57226 => x"10",		-- 00df8a: 104B             BR      0x0014(R11)
						   57227 => x"6B",
						   57228 => x"14",		-- 00df8c: 1400            
						   57229 => x"00",
						   57230 => x"3C",		-- 00df8e: 3C43             MOV.W   #-1,R12
						   57231 => x"63",
						   57232 => x"3D",		-- 00df90: 3D43             MOV.W   #-1,R13
						   57233 => x"63",
						   57234 => x"30",		-- 00df92: 3041             RET     
						   57235 => x"61",
						   -- Begin: __mspabi_mpyl
						   -- Begin: __mspabi_mpyl_sw
						   57236 => x"0A",		-- 00df94: 0A12             PUSH    R10
						   57237 => x"32",
						   57238 => x"0A",		-- 00df96: 0A43             CLR.W   R10
						   57239 => x"63",
						   57240 => x"0B",		-- 00df98: 0B43             CLR.W   R11
						   57241 => x"63",
						   -- Begin: mpyl_add_loop
						   57242 => x"12",		-- 00df9a: 12C3             CLRC    
						   57243 => x"E3",
						   57244 => x"0D",		-- 00df9c: 0D10             RRC     R13
						   57245 => x"30",
						   57246 => x"0C",		-- 00df9e: 0C10             RRC     R12
						   57247 => x"30",
						   57248 => x"02",		-- 00dfa0: 0228             JLO     (shift_test_mpyl)
						   57249 => x"48",
						   57250 => x"0A",		-- 00dfa2: 0A5E             ADD.W   R14,R10
						   57251 => x"7E",
						   57252 => x"0B",		-- 00dfa4: 0B6F             ADDC.W  R15,R11
						   57253 => x"8F",
						   -- Begin: shift_test_mpyl
						   57254 => x"0E",		-- 00dfa6: 0E5E             RLA.W   R14
						   57255 => x"7E",
						   57256 => x"0F",		-- 00dfa8: 0F6F             RLC.W   R15
						   57257 => x"8F",
						   57258 => x"0D",		-- 00dfaa: 0D93             TST.W   R13
						   57259 => x"B3",
						   57260 => x"F6",		-- 00dfac: F623             JNE     (mpyl_add_loop)
						   57261 => x"43",
						   57262 => x"0C",		-- 00dfae: 0C93             TST.W   R12
						   57263 => x"B3",
						   57264 => x"F4",		-- 00dfb0: F423             JNE     (mpyl_add_loop)
						   57265 => x"43",
						   57266 => x"0C",		-- 00dfb2: 0C4A             MOV.W   R10,R12
						   57267 => x"6A",
						   57268 => x"0D",		-- 00dfb4: 0D4B             MOV.W   R11,R13
						   57269 => x"6B",
						   57270 => x"3A",		-- 00dfb6: 3A41             POP.W   R10
						   57271 => x"61",
						   57272 => x"30",		-- 00dfb8: 3041             RET     
						   57273 => x"61",
						   -- Begin: write
						   57274 => x"0C",		-- 00dfba: 0C93             TST.W   R12
						   57275 => x"B3",
						   57276 => x"0E",		-- 00dfbc: 0E38             JL      ($C$L1)
						   57277 => x"58",
						   57278 => x"3C",		-- 00dfbe: 3C90             CMP.W   #0x000a,R12
						   57279 => x"B0",
						   57280 => x"0A",		-- 00dfc0: 0A00            
						   57281 => x"00",
						   57282 => x"0B",		-- 00dfc2: 0B34             JGE     ($C$L1)
						   57283 => x"54",
						   57284 => x"0C",		-- 00dfc4: 0C5C             RLA.W   R12
						   57285 => x"7C",
						   57286 => x"0C",		-- 00dfc6: 0C5C             RLA.W   R12
						   57287 => x"7C",
						   57288 => x"3C",		-- 00dfc8: 3C50             ADD.W   #0x20c6,R12
						   57289 => x"70",
						   57290 => x"C6",		-- 00dfca: C620            
						   57291 => x"20",
						   57292 => x"2F",		-- 00dfcc: 2F4C             MOV.W   @R12,R15
						   57293 => x"6C",
						   57294 => x"0F",		-- 00dfce: 0F93             TST.W   R15
						   57295 => x"B3",
						   57296 => x"04",		-- 00dfd0: 0424             JEQ     ($C$L1)
						   57297 => x"44",
						   57298 => x"1C",		-- 00dfd2: 1C4C             MOV.W   0x0002(R12),R12
						   57299 => x"6C",
						   57300 => x"02",		-- 00dfd4: 0200            
						   57301 => x"00",
						   57302 => x"10",		-- 00dfd6: 104F             BR      0x0012(R15)
						   57303 => x"6F",
						   57304 => x"12",		-- 00dfd8: 1200            
						   57305 => x"00",
						   57306 => x"3C",		-- 00dfda: 3C43             MOV.W   #-1,R12
						   57307 => x"63",
						   57308 => x"30",		-- 00dfdc: 3041             RET     
						   57309 => x"61",
						   -- Begin: __mspabi_mpyul
						   -- Begin: __mspabi_mpyul_sw
						   57310 => x"0B",		-- 00dfde: 0B4C             MOV.W   R12,R11
						   57311 => x"6C",
						   57312 => x"0E",		-- 00dfe0: 0E4D             MOV.W   R13,R14
						   57313 => x"6D",
						   57314 => x"0F",		-- 00dfe2: 0F43             CLR.W   R15
						   57315 => x"63",
						   57316 => x"0C",		-- 00dfe4: 0C43             CLR.W   R12
						   57317 => x"63",
						   57318 => x"0D",		-- 00dfe6: 0D43             CLR.W   R13
						   57319 => x"63",
						   57320 => x"12",		-- 00dfe8: 12C3             CLRC    
						   57321 => x"E3",
						   57322 => x"0B",		-- 00dfea: 0B10             RRC     R11
						   57323 => x"30",
						   57324 => x"01",		-- 00dfec: 013C             JMP     (mpyul_add_loop1)
						   57325 => x"5C",
						   -- Begin: mpyul_add_loop
						   57326 => x"0B",		-- 00dfee: 0B11             RRA     R11
						   57327 => x"31",
						   -- Begin: mpyul_add_loop1
						   57328 => x"02",		-- 00dff0: 0228             JLO     (shift_test_mpyul)
						   57329 => x"48",
						   57330 => x"0C",		-- 00dff2: 0C5E             ADD.W   R14,R12
						   57331 => x"7E",
						   57332 => x"0D",		-- 00dff4: 0D6F             ADDC.W  R15,R13
						   57333 => x"8F",
						   -- Begin: shift_test_mpyul
						   57334 => x"0E",		-- 00dff6: 0E5E             RLA.W   R14
						   57335 => x"7E",
						   57336 => x"0F",		-- 00dff8: 0F6F             RLC.W   R15
						   57337 => x"8F",
						   57338 => x"0B",		-- 00dffa: 0B93             TST.W   R11
						   57339 => x"B3",
						   57340 => x"F8",		-- 00dffc: F823             JNE     (mpyul_add_loop)
						   57341 => x"43",
						   57342 => x"30",		-- 00dffe: 3041             RET     
						   57343 => x"61",
						   -- Begin: memccpy
						   57344 => x"0A",		-- 00e000: 0A12             PUSH    R10
						   57345 => x"32",
						   57346 => x"0F",		-- 00e002: 0F93             TST.W   R15
						   57347 => x"B3",
						   57348 => x"0B",		-- 00e004: 0B24             JEQ     ($C$L2)
						   57349 => x"44",
						   57350 => x"4E",		-- 00e006: 4E4E             MOV.B   R14,R14
						   57351 => x"6E",
						   57352 => x"6B",		-- 00e008: 6B4D             MOV.B   @R13,R11
						   57353 => x"6D",
						   57354 => x"1C",		-- 00e00a: 1C53             INC.W   R12
						   57355 => x"73",
						   57356 => x"CC",		-- 00e00c: CC4B             MOV.B   R11,0xffff(R12)
						   57357 => x"6B",
						   57358 => x"FF",		-- 00e00e: FFFF            
						   57359 => x"FF",
						   57360 => x"4A",		-- 00e010: 4A4E             MOV.B   R14,R10
						   57361 => x"6E",
						   57362 => x"0B",		-- 00e012: 0B9A             CMP.W   R10,R11
						   57363 => x"BA",
						   57364 => x"04",		-- 00e014: 0424             JEQ     ($C$L3)
						   57365 => x"44",
						   57366 => x"1D",		-- 00e016: 1D53             INC.W   R13
						   57367 => x"73",
						   57368 => x"1F",		-- 00e018: 1F83             DEC.W   R15
						   57369 => x"A3",
						   57370 => x"F6",		-- 00e01a: F623             JNE     ($C$L1)
						   57371 => x"43",
						   57372 => x"0C",		-- 00e01c: 0C43             CLR.W   R12
						   57373 => x"63",
						   57374 => x"3A",		-- 00e01e: 3A41             POP.W   R10
						   57375 => x"61",
						   57376 => x"30",		-- 00e020: 3041             RET     
						   57377 => x"61",
						   -- Begin: __mspabi_mpyull
						   -- Begin: __mspabi_mpyull_sw
						   57378 => x"0A",		-- 00e022: 0A12             PUSH    R10
						   57379 => x"32",
						   57380 => x"09",		-- 00e024: 0912             PUSH    R9
						   57381 => x"32",
						   57382 => x"08",		-- 00e026: 0812             PUSH    R8
						   57383 => x"32",
						   57384 => x"08",		-- 00e028: 084C             MOV.W   R12,R8
						   57385 => x"6C",
						   57386 => x"09",		-- 00e02a: 094D             MOV.W   R13,R9
						   57387 => x"6D",
						   57388 => x"0A",		-- 00e02c: 0A43             CLR.W   R10
						   57389 => x"63",
						   57390 => x"0B",		-- 00e02e: 0B43             CLR.W   R11
						   57391 => x"63",
						   57392 => x"0C",		-- 00e030: 0C4E             MOV.W   R14,R12
						   57393 => x"6E",
						   57394 => x"0D",		-- 00e032: 0D4F             MOV.W   R15,R13
						   57395 => x"6F",
						   57396 => x"0E",		-- 00e034: 0E43             CLR.W   R14
						   57397 => x"63",
						   57398 => x"0F",		-- 00e036: 0F43             CLR.W   R15
						   57399 => x"63",
						   57400 => x"B0",		-- 00e038: B012             CALL    #__mspabi_mpyll_sw
						   57401 => x"32",
						   57402 => x"D6",		-- 00e03a: D6C5            
						   57403 => x"C5",
						   57404 => x"30",		-- 00e03c: 3040             BR      #__mspabi_func_epilog_3
						   57405 => x"60",
						   57406 => x"62",		-- 00e03e: 62E1            
						   57407 => x"E1",
						   -- Begin: _c_int00_noargs
						   57408 => x"31",		-- 00e040: 3140             MOV.W   #0x3000,SP
						   57409 => x"60",
						   57410 => x"00",		-- 00e042: 0030            
						   57411 => x"30",
						   57412 => x"B0",		-- 00e044: B012             CALL    #_system_pre_init
						   57413 => x"32",
						   57414 => x"C2",		-- 00e046: C2E1            
						   57415 => x"E1",
						   57416 => x"0C",		-- 00e048: 0C93             TST.W   R12
						   57417 => x"B3",
						   57418 => x"02",		-- 00e04a: 0224             JEQ     ($C$L2)
						   57419 => x"44",
						   57420 => x"B0",		-- 00e04c: B012             CALL    #__TI_auto_init_nobinit_nopinit
						   57421 => x"32",
						   57422 => x"B0",		-- 00e04e: B0DB            
						   57423 => x"DB",
						   57424 => x"0C",		-- 00e050: 0C43             CLR.W   R12
						   57425 => x"63",
						   57426 => x"B0",		-- 00e052: B012             CALL    #main
						   57427 => x"32",
						   57428 => x"54",		-- 00e054: 54DA            
						   57429 => x"DA",
						   57430 => x"1C",		-- 00e056: 1C43             MOV.W   #1,R12
						   57431 => x"63",
						   57432 => x"B0",		-- 00e058: B012             CALL    #exit
						   57433 => x"32",
						   57434 => x"6C",		-- 00e05a: 6CDB            
						   57435 => x"DB",
						   -- Begin: free_list_remove
						   57436 => x"3F",		-- 00e05c: 3F40             MOV.W   #0x21a6,R15
						   57437 => x"60",
						   57438 => x"A6",		-- 00e05e: A621            
						   57439 => x"21",
						   57440 => x"02",		-- 00e060: 023C             JMP     ($C$L2)
						   57441 => x"5C",
						   57442 => x"2F",		-- 00e062: 2F42             MOV.W   #4,R15
						   57443 => x"62",
						   57444 => x"0F",		-- 00e064: 0F5E             ADD.W   R14,R15
						   57445 => x"7E",
						   57446 => x"2E",		-- 00e066: 2E4F             MOV.W   @R15,R14
						   57447 => x"6F",
						   57448 => x"0E",		-- 00e068: 0E93             TST.W   R14
						   57449 => x"B3",
						   57450 => x"05",		-- 00e06a: 0524             JEQ     ($C$L3)
						   57451 => x"44",
						   57452 => x"0E",		-- 00e06c: 0E9C             CMP.W   R12,R14
						   57453 => x"BC",
						   57454 => x"F9",		-- 00e06e: F923             JNE     ($C$L1)
						   57455 => x"43",
						   57456 => x"9F",		-- 00e070: 9F4C             MOV.W   0x0004(R12),0x0000(R15)
						   57457 => x"6C",
						   57458 => x"04",		-- 00e072: 0400            
						   57459 => x"00",
						   57460 => x"00",		-- 00e074: 0000            
						   57461 => x"00",
						   57462 => x"30",		-- 00e076: 3041             RET     
						   57463 => x"61",
						   -- Begin: strchr
						   57464 => x"6F",		-- 00e078: 6F4C             MOV.B   @R12,R15
						   57465 => x"6C",
						   57466 => x"4D",		-- 00e07a: 4D4D             MOV.B   R13,R13
						   57467 => x"6D",
						   57468 => x"06",		-- 00e07c: 063C             JMP     ($C$L3)
						   57469 => x"5C",
						   57470 => x"0F",		-- 00e07e: 0F93             TST.W   R15
						   57471 => x"B3",
						   57472 => x"02",		-- 00e080: 0220             JNE     ($C$L2)
						   57473 => x"40",
						   57474 => x"0C",		-- 00e082: 0C43             CLR.W   R12
						   57475 => x"63",
						   57476 => x"30",		-- 00e084: 3041             RET     
						   57477 => x"61",
						   57478 => x"1C",		-- 00e086: 1C53             INC.W   R12
						   57479 => x"73",
						   57480 => x"6F",		-- 00e088: 6F4C             MOV.B   @R12,R15
						   57481 => x"6C",
						   57482 => x"4E",		-- 00e08a: 4E4D             MOV.B   R13,R14
						   57483 => x"6D",
						   57484 => x"0F",		-- 00e08c: 0F9E             CMP.W   R14,R15
						   57485 => x"BE",
						   57486 => x"F7",		-- 00e08e: F723             JNE     ($C$L1)
						   57487 => x"43",
						   57488 => x"30",		-- 00e090: 3041             RET     
						   57489 => x"61",
						   -- Begin: strcmp
						   57490 => x"0F",		-- 00e092: 0F4C             MOV.W   R12,R15
						   57491 => x"6C",
						   57492 => x"6E",		-- 00e094: 6E4F             MOV.B   @R15,R14
						   57493 => x"6F",
						   57494 => x"6B",		-- 00e096: 6B4D             MOV.B   @R13,R11
						   57495 => x"6D",
						   57496 => x"4C",		-- 00e098: 4C4E             MOV.B   R14,R12
						   57497 => x"6E",
						   57498 => x"0C",		-- 00e09a: 0C8B             SUB.W   R11,R12
						   57499 => x"AB",
						   57500 => x"4E",		-- 00e09c: 4E93             TST.B   R14
						   57501 => x"B3",
						   57502 => x"04",		-- 00e09e: 0424             JEQ     ($C$L2)
						   57503 => x"44",
						   57504 => x"1D",		-- 00e0a0: 1D53             INC.W   R13
						   57505 => x"73",
						   57506 => x"1F",		-- 00e0a2: 1F53             INC.W   R15
						   57507 => x"73",
						   57508 => x"0C",		-- 00e0a4: 0C93             TST.W   R12
						   57509 => x"B3",
						   57510 => x"F6",		-- 00e0a6: F627             JEQ     ($C$L1)
						   57511 => x"47",
						   57512 => x"30",		-- 00e0a8: 3041             RET     
						   57513 => x"61",
						   -- Begin: __mspabi_divu
						   -- Begin: __mspabi_remu
						   57514 => x"0E",		-- 00e0aa: 0E43             CLR.W   R14
						   57515 => x"63",
						   57516 => x"0F",		-- 00e0ac: 0F4C             MOV.W   R12,R15
						   57517 => x"6C",
						   57518 => x"1C",		-- 00e0ae: 1C43             MOV.W   #1,R12
						   57519 => x"63",
						   -- Begin: div_loop
						   57520 => x"0F",		-- 00e0b0: 0F5F             RLA.W   R15
						   57521 => x"7F",
						   57522 => x"0E",		-- 00e0b2: 0E6E             RLC.W   R14
						   57523 => x"8E",
						   57524 => x"0E",		-- 00e0b4: 0E9D             CMP.W   R13,R14
						   57525 => x"BD",
						   57526 => x"01",		-- 00e0b6: 0128             JLO     (set_quotient_bit)
						   57527 => x"48",
						   57528 => x"0E",		-- 00e0b8: 0E8D             SUB.W   R13,R14
						   57529 => x"AD",
						   -- Begin: set_quotient_bit
						   57530 => x"0C",		-- 00e0ba: 0C6C             RLC.W   R12
						   57531 => x"8C",
						   57532 => x"F9",		-- 00e0bc: F92B             JLO     (div_loop)
						   57533 => x"4B",
						   57534 => x"30",		-- 00e0be: 3041             RET     
						   57535 => x"61",
						   -- Begin: __TI_zero_init_nomemset
						   57536 => x"1F",		-- 00e0c0: 1F4C             MOV.W   0x0001(R12),R15
						   57537 => x"6C",
						   57538 => x"01",		-- 00e0c2: 0100            
						   57539 => x"00",
						   57540 => x"0F",		-- 00e0c4: 0F93             TST.W   R15
						   57541 => x"B3",
						   57542 => x"05",		-- 00e0c6: 0524             JEQ     ($C$L2)
						   57543 => x"44",
						   57544 => x"1D",		-- 00e0c8: 1D53             INC.W   R13
						   57545 => x"73",
						   57546 => x"CD",		-- 00e0ca: CD43             CLR.B   0xffff(R13)
						   57547 => x"63",
						   57548 => x"FF",		-- 00e0cc: FFFF            
						   57549 => x"FF",
						   57550 => x"1F",		-- 00e0ce: 1F83             DEC.W   R15
						   57551 => x"A3",
						   57552 => x"FB",		-- 00e0d0: FB23             JNE     ($C$L1)
						   57553 => x"43",
						   57554 => x"30",		-- 00e0d2: 3041             RET     
						   57555 => x"61",
						   -- Begin: memchr
						   57556 => x"0E",		-- 00e0d4: 0E93             TST.W   R14
						   57557 => x"B3",
						   57558 => x"06",		-- 00e0d6: 0624             JEQ     ($C$L2)
						   57559 => x"44",
						   57560 => x"4D",		-- 00e0d8: 4D4D             MOV.B   R13,R13
						   57561 => x"6D",
						   57562 => x"6D",		-- 00e0da: 6D9C             CMP.B   @R12,R13
						   57563 => x"BC",
						   57564 => x"04",		-- 00e0dc: 0424             JEQ     ($C$L3)
						   57565 => x"44",
						   57566 => x"1C",		-- 00e0de: 1C53             INC.W   R12
						   57567 => x"73",
						   57568 => x"1E",		-- 00e0e0: 1E83             DEC.W   R14
						   57569 => x"A3",
						   57570 => x"FB",		-- 00e0e2: FB23             JNE     ($C$L1)
						   57571 => x"43",
						   57572 => x"0C",		-- 00e0e4: 0C43             CLR.W   R12
						   57573 => x"63",
						   57574 => x"30",		-- 00e0e6: 3041             RET     
						   57575 => x"61",
						   -- Begin: memset
						   57576 => x"0F",		-- 00e0e8: 0F4C             MOV.W   R12,R15
						   57577 => x"6C",
						   57578 => x"0E",		-- 00e0ea: 0E93             TST.W   R14
						   57579 => x"B3",
						   57580 => x"06",		-- 00e0ec: 0624             JEQ     ($C$L2)
						   57581 => x"44",
						   57582 => x"4D",		-- 00e0ee: 4D4D             MOV.B   R13,R13
						   57583 => x"6D",
						   57584 => x"1F",		-- 00e0f0: 1F53             INC.W   R15
						   57585 => x"73",
						   57586 => x"CF",		-- 00e0f2: CF4D             MOV.B   R13,0xffff(R15)
						   57587 => x"6D",
						   57588 => x"FF",		-- 00e0f4: FFFF            
						   57589 => x"FF",
						   57590 => x"1E",		-- 00e0f6: 1E83             DEC.W   R14
						   57591 => x"A3",
						   57592 => x"FB",		-- 00e0f8: FB23             JNE     ($C$L1)
						   57593 => x"43",
						   57594 => x"30",		-- 00e0fa: 3041             RET     
						   57595 => x"61",
						   -- Begin: __mspabi_mpyi
						   -- Begin: __mspabi_mpyi_sw
						   57596 => x"0E",		-- 00e0fc: 0E43             CLR.W   R14
						   57597 => x"63",
						   -- Begin: mpyi_add_loop
						   57598 => x"12",		-- 00e0fe: 12C3             CLRC    
						   57599 => x"E3",
						   57600 => x"0C",		-- 00e100: 0C10             RRC     R12
						   57601 => x"30",
						   57602 => x"01",		-- 00e102: 0128             JLO     (shift_test_mpyi)
						   57603 => x"48",
						   57604 => x"0E",		-- 00e104: 0E5D             ADD.W   R13,R14
						   57605 => x"7D",
						   -- Begin: shift_test_mpyi
						   57606 => x"0D",		-- 00e106: 0D5D             RLA.W   R13
						   57607 => x"7D",
						   57608 => x"0C",		-- 00e108: 0C93             TST.W   R12
						   57609 => x"B3",
						   57610 => x"F9",		-- 00e10a: F923             JNE     (mpyi_add_loop)
						   57611 => x"43",
						   57612 => x"0C",		-- 00e10c: 0C4E             MOV.W   R14,R12
						   57613 => x"6E",
						   57614 => x"30",		-- 00e10e: 3041             RET     
						   57615 => x"61",
						   -- Begin: wcslen
						   57616 => x"0F",		-- 00e110: 0F4C             MOV.W   R12,R15
						   57617 => x"6C",
						   57618 => x"01",		-- 00e112: 013C             JMP     ($C$L2)
						   57619 => x"5C",
						   57620 => x"2F",		-- 00e114: 2F53             INCD.W  R15
						   57621 => x"73",
						   57622 => x"8F",		-- 00e116: 8F93             TST.W   0x0000(R15)
						   57623 => x"B3",
						   57624 => x"00",		-- 00e118: 0000            
						   57625 => x"00",
						   57626 => x"FC",		-- 00e11a: FC23             JNE     ($C$L1)
						   57627 => x"43",
						   57628 => x"0F",		-- 00e11c: 0F8C             SUB.W   R12,R15
						   57629 => x"AC",
						   57630 => x"0F",		-- 00e11e: 0F11             RRA     R15
						   57631 => x"31",
						   57632 => x"0C",		-- 00e120: 0C4F             MOV.W   R15,R12
						   57633 => x"6F",
						   57634 => x"30",		-- 00e122: 3041             RET     
						   57635 => x"61",
						   -- Begin: __TI_decompress_none
						   57636 => x"0F",		-- 00e124: 0F4C             MOV.W   R12,R15
						   57637 => x"6C",
						   57638 => x"0C",		-- 00e126: 0C4D             MOV.W   R13,R12
						   57639 => x"6D",
						   57640 => x"3D",		-- 00e128: 3D40             MOV.W   #0x0003,R13
						   57641 => x"60",
						   57642 => x"03",		-- 00e12a: 0300            
						   57643 => x"00",
						   57644 => x"0D",		-- 00e12c: 0D5F             ADD.W   R15,R13
						   57645 => x"7F",
						   57646 => x"1E",		-- 00e12e: 1E4F             MOV.W   0x0001(R15),R14
						   57647 => x"6F",
						   57648 => x"01",		-- 00e130: 0100            
						   57649 => x"00",
						   57650 => x"30",		-- 00e132: 3040             BR      #memcpy
						   57651 => x"60",
						   57652 => x"48",		-- 00e134: 48E1            
						   57653 => x"E1",
						   -- Begin: __mspabi_srll
						   57654 => x"3E",		-- 00e136: 3EF0             AND.W   #0x001f,R14
						   57655 => x"10",
						   57656 => x"1F",		-- 00e138: 1F00            
						   57657 => x"00",
						   57658 => x"05",		-- 00e13a: 0524             JEQ     (L_LSR_RET)
						   57659 => x"44",
						   -- Begin: L_LSR_TOP
						   57660 => x"12",		-- 00e13c: 12C3             CLRC    
						   57661 => x"E3",
						   57662 => x"0D",		-- 00e13e: 0D10             RRC     R13
						   57663 => x"30",
						   57664 => x"0C",		-- 00e140: 0C10             RRC     R12
						   57665 => x"30",
						   57666 => x"1E",		-- 00e142: 1E83             DEC.W   R14
						   57667 => x"A3",
						   57668 => x"FB",		-- 00e144: FB23             JNE     (L_LSR_TOP)
						   57669 => x"43",
						   -- Begin: L_LSR_RET
						   57670 => x"30",		-- 00e146: 3041             RET     
						   57671 => x"61",
						   -- Begin: memcpy
						   57672 => x"0E",		-- 00e148: 0E93             TST.W   R14
						   57673 => x"B3",
						   57674 => x"06",		-- 00e14a: 0624             JEQ     ($C$L2)
						   57675 => x"44",
						   57676 => x"0F",		-- 00e14c: 0F4C             MOV.W   R12,R15
						   57677 => x"6C",
						   57678 => x"1F",		-- 00e14e: 1F53             INC.W   R15
						   57679 => x"73",
						   57680 => x"FF",		-- 00e150: FF4D             MOV.B   @R13+,0xffff(R15)
						   57681 => x"6D",
						   57682 => x"FF",		-- 00e152: FFFF            
						   57683 => x"FF",
						   57684 => x"1E",		-- 00e154: 1E83             DEC.W   R14
						   57685 => x"A3",
						   57686 => x"FB",		-- 00e156: FB23             JNE     ($C$L1)
						   57687 => x"43",
						   57688 => x"30",		-- 00e158: 3041             RET     
						   57689 => x"61",
						   -- Begin: __mspabi_func_epilog_7
						   -- Begin: __mspabi_func_epilog
						   57690 => x"34",		-- 00e15a: 3441             POP.W   R4
						   57691 => x"61",
						   -- Begin: __mspabi_func_epilog_6
						   57692 => x"35",		-- 00e15c: 3541             POP.W   R5
						   57693 => x"61",
						   -- Begin: __mspabi_func_epilog_5
						   57694 => x"36",		-- 00e15e: 3641             POP.W   R6
						   57695 => x"61",
						   -- Begin: __mspabi_func_epilog_4
						   57696 => x"37",		-- 00e160: 3741             POP.W   R7
						   57697 => x"61",
						   -- Begin: __mspabi_func_epilog_3
						   57698 => x"38",		-- 00e162: 3841             POP.W   R8
						   57699 => x"61",
						   -- Begin: __mspabi_func_epilog_2
						   57700 => x"39",		-- 00e164: 3941             POP.W   R9
						   57701 => x"61",
						   -- Begin: __mspabi_func_epilog_1
						   57702 => x"3A",		-- 00e166: 3A41             POP.W   R10
						   57703 => x"61",
						   57704 => x"30",		-- 00e168: 3041             RET     
						   57705 => x"61",
						   -- Begin: strcpy
						   57706 => x"0F",		-- 00e16a: 0F4C             MOV.W   R12,R15
						   57707 => x"6C",
						   57708 => x"7E",		-- 00e16c: 7E4D             MOV.B   @R13+,R14
						   57709 => x"6D",
						   57710 => x"1F",		-- 00e16e: 1F53             INC.W   R15
						   57711 => x"73",
						   57712 => x"CF",		-- 00e170: CF4E             MOV.B   R14,0xffff(R15)
						   57713 => x"6E",
						   57714 => x"FF",		-- 00e172: FFFF            
						   57715 => x"FF",
						   57716 => x"0E",		-- 00e174: 0E93             TST.W   R14
						   57717 => x"B3",
						   57718 => x"FA",		-- 00e176: FA23             JNE     ($C$L1)
						   57719 => x"43",
						   57720 => x"30",		-- 00e178: 3041             RET     
						   57721 => x"61",
						   -- Begin: strlen
						   57722 => x"3F",		-- 00e17a: 3F43             MOV.W   #-1,R15
						   57723 => x"63",
						   57724 => x"1F",		-- 00e17c: 1F53             INC.W   R15
						   57725 => x"73",
						   57726 => x"7E",		-- 00e17e: 7E4C             MOV.B   @R12+,R14
						   57727 => x"6C",
						   57728 => x"0E",		-- 00e180: 0E93             TST.W   R14
						   57729 => x"B3",
						   57730 => x"FC",		-- 00e182: FC23             JNE     ($C$L1)
						   57731 => x"43",
						   57732 => x"0C",		-- 00e184: 0C4F             MOV.W   R15,R12
						   57733 => x"6F",
						   57734 => x"30",		-- 00e186: 3041             RET     
						   57735 => x"61",
						   -- Begin: __mspabi_fltid
						   57736 => x"3C",		-- 00e188: 3CB0             BIT.W   #0x8000,R12
						   57737 => x"D0",
						   57738 => x"00",		-- 00e18a: 0080            
						   57739 => x"80",
						   57740 => x"0D",		-- 00e18c: 0D7D             SUBC.W  R13,R13
						   57741 => x"9D",
						   57742 => x"3D",		-- 00e18e: 3DE3             INV.W   R13
						   57743 => x"03",
						   57744 => x"30",		-- 00e190: 3040             BR      #__mspabi_fltlid
						   57745 => x"60",
						   57746 => x"94",		-- 00e192: 94CE            
						   57747 => x"CE",
						   -- Begin: toupper
						   57748 => x"EC",		-- 00e194: ECB3             BIT.B   #2,0x9917(R12)
						   57749 => x"D3",
						   57750 => x"17",		-- 00e196: 1799            
						   57751 => x"99",
						   57752 => x"02",		-- 00e198: 0224             JEQ     ($C$L1)
						   57753 => x"44",
						   57754 => x"3C",		-- 00e19a: 3C80             SUB.W   #0x0020,R12
						   57755 => x"A0",
						   57756 => x"20",		-- 00e19c: 2000            
						   57757 => x"00",
						   57758 => x"30",		-- 00e19e: 3041             RET     
						   57759 => x"61",
						   -- Begin: abs
						   57760 => x"0C",		-- 00e1a0: 0C93             TST.W   R12
						   57761 => x"B3",
						   57762 => x"02",		-- 00e1a2: 0234             JGE     ($C$L1)
						   57763 => x"54",
						   57764 => x"3C",		-- 00e1a4: 3CE3             INV.W   R12
						   57765 => x"03",
						   57766 => x"1C",		-- 00e1a6: 1C53             INC.W   R12
						   57767 => x"73",
						   57768 => x"30",		-- 00e1a8: 3041             RET     
						   57769 => x"61",
						   -- Begin: malloc
						   57770 => x"0D",		-- 00e1aa: 0D4C             MOV.W   R12,R13
						   57771 => x"6C",
						   57772 => x"2C",		-- 00e1ac: 2C42             MOV.W   #4,R12
						   57773 => x"62",
						   57774 => x"30",		-- 00e1ae: 3040             BR      #aligned_alloc
						   57775 => x"60",
						   57776 => x"E2",		-- 00e1b0: E2C7            
						   57777 => x"C7",
						   -- Begin: _outc
						   57778 => x"4C",		-- 00e1b2: 4C4C             MOV.B   R12,R12
						   57779 => x"6C",
						   57780 => x"30",		-- 00e1b4: 3040             BR      #fputc
						   57781 => x"60",
						   57782 => x"7E",		-- 00e1b6: 7ED0            
						   57783 => x"D0",
						   -- Begin: abort
						   57784 => x"03",		-- 00e1b8: 0343             NOP     
						   57785 => x"63",
						   57786 => x"FF",		-- 00e1ba: FF3F             JMP     ($C$L1)
						   57787 => x"5F",
						   57788 => x"03",		-- 00e1bc: 0343             NOP     
						   57789 => x"63",
						   -- Begin: _outs
						   57790 => x"30",		-- 00e1be: 3040             BR      #fputs
						   57791 => x"60",
						   57792 => x"D8",		-- 00e1c0: D8C8            
						   57793 => x"C8",
						   -- Begin: _system_pre_init
						   57794 => x"1C",		-- 00e1c2: 1C43             MOV.W   #1,R12
						   57795 => x"63",
						   57796 => x"30",		-- 00e1c4: 3041             RET     
						   57797 => x"61",
						   -- Begin: _nop
						   57798 => x"30",		-- 00e1c6: 3041             RET     
						   57799 => x"61",
						   -- Begin: _system_post_cinit
						   57800 => x"30",		-- 00e1c8: 3041             RET     
						   57801 => x"61",
						   -- ISR Trap
						   57802 => x"32",		-- 00e1ca: 32D0             BIS.W   #0x0010,SR
						   57803 => x"F0",
						   57804 => x"10",		-- 00e1cc: 1000            
						   57805 => x"00",
						   57806 => x"FD",		-- 00e1ce: FD3F             JMP     (__TI_ISR_TRAP)
						   57807 => x"5F",
						   57808 => x"03",		-- 00e1d0: 0343             NOP     
						   57809 => x"63",
						   -- IRQ Vectors (Interrupt Vectors)
						   65486 => x"ca",		-- 00ffce:e1ca PORT4 __TI_int22 int22
						   65487 => x"e1",
						   65488 => x"ca",		-- 00ffd0:e1ca PORT3 __TI_int23 int23
						   65489 => x"e1",
						   65490 => x"ca",		-- 00ffd2:e1ca PORT2 __TI_int24 int24
						   65491 => x"e1",
						   65492 => x"ca",		-- 00ffd4:e1ca PORT1 __TI_int25 int25
						   65493 => x"e1",
						   65494 => x"ca",		-- 00ffd6:e1ca SAC1_SAC3 __TI_int26 int26
						   65495 => x"e1",
						   65496 => x"ca",		-- 00ffd8:e1ca SAC0_SAC2 __TI_int27 int27
						   65497 => x"e1",
						   65498 => x"ca",		-- 00ffda:e1ca ECOMP0_ECOMP1 __TI_int28 int28
						   65499 => x"e1",
						   65500 => x"ca",		-- 00ffdc:e1ca ADC __TI_int29 int29
						   65501 => x"e1",
						   65502 => x"ca",		-- 00ffde:e1ca EUSCI_B1 __TI_int30 int30
						   65503 => x"e1",
						   65504 => x"ca",		-- 00ffe0:e1ca EUSCI_B0 __TI_int31 int31
						   65505 => x"e1",
						   65506 => x"ca",		-- 00ffe2:e1ca EUSCI_A1 __TI_int32 int32
						   65507 => x"e1",
						   65508 => x"ca",		-- 00ffe4:e1ca EUSCI_A0 __TI_int33 int33
						   65509 => x"e1",
						   65510 => x"ca",		-- 00ffe6:e1ca WDT __TI_int34 int34
						   65511 => x"e1",
						   65512 => x"ca",		-- 00ffe8:e1ca RTC __TI_int35 int35
						   65513 => x"e1",
						   65514 => x"ca",		-- 00ffea:e1ca TIMER3_B1 __TI_int36 int36
						   65515 => x"e1",
						   65516 => x"ca",		-- 00ffec:e1ca TIMER3_B0 __TI_int37 int37
						   65517 => x"e1",
						   65518 => x"ca",		-- 00ffee:e1ca TIMER2_B1 __TI_int38 int38
						   65519 => x"e1",
						   65520 => x"ca",		-- 00fff0:e1ca TIMER2_B0 __TI_int39 int39
						   65521 => x"e1",
						   65522 => x"ca",		-- 00fff2:e1ca TIMER1_B1 __TI_int40 int40
						   65523 => x"e1",
						   65524 => x"ca",		-- 00fff4:e1ca TIMER1_B0 __TI_int41 int41
						   65525 => x"e1",
						   65526 => x"ca",		-- 00fff6:e1ca TIMER0_B1 __TI_int42 int42
						   65527 => x"e1",
						   65528 => x"ca",		-- 00fff8:e1ca TIMER0_B0 __TI_int43 int43
						   65529 => x"e1",
						   65530 => x"ca",		-- 00fffa:e1ca UNMI __TI_int44 int44
						   65531 => x"e1",
						   65532 => x"ca",		-- 00fffc:e1ca SYSNMI __TI_int45 int45
						   65533 => x"e1",

                           65534 =>  x"00",		-- Reset Vector = xFFFE:xFFFF
                           65535 =>  x"80",		--  Startup Value = x8000

                           others => x"00");

    signal EN : std_logic;
    
    begin
    -- Note 1:  The bus system uses a 16-bit Address (MAB)
    --          This address size can access locations from x0000 to xFFFF
    --          But our array is only defined from x8000 to xFFFF and
    --          if we try to access it with any other address, it will crash.
    --          So the first thing we need to do is create a local enable that
    --          will only assert when MAB is within x8000 to xFFFF.

     LOCAL_EN : process (MAB) 
     begin
         if ( (to_integer(unsigned(MAB)) >= 32768) and (to_integer(unsigned(MAB)) <= 65535)) then
           EN <= '1';
         else 
           EN <= '0';
         end if;
     end process;

    
    -- Note 2:  The bus system uses a 16-bit Address (MAB)
    --          The MDB_out is also provided as a 16-bit word
    --          However, the memory array is actually built as 8-bit bytes.
    --          So for a given 16-bit MAB, we give MDB_out = HB : LB
    --                                                 or  = ROM(MAB);1) : ROM(MAB)

    MEMORY_ROM : process (clk) 
    begin
        if (rising_edge(clk)) then
            if (EN='1' and write='0') then                      
              MDB_in <= ROM(to_integer(unsigned(MAB)) + 1 ) & ROM(to_integer(unsigned(MAB))); 
            end if;
        end if;
    end process;


end architecture;