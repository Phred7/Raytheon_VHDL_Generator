library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;


entity highroller_memory is
    port ( clk	: in	std_logic;
         MAB		: in	std_logic_vector(15 downto 0);
         MDB_in  	: out	std_logic_vector(15 downto 0);
         MDB_out  	: in	std_logic_vector(15 downto 0);
         write	    : in	std_logic);
end entity;

architecture highroller_memory_arch of highroller_memory is

type rom_type is array (32768 to 65535) of std_logic_vector(7 downto 0);  -- this is MAB: x8000 to xFFFF
    
constant ROM : rom_type :=(32768 => x"31",		-- 008000: 3140             MOV.W   #0x3000,SP
						   32769 => x"60",
						   32770 => x"00",		-- 008002: 0030            
						   32771 => x"30",
						   32772 => x"B2",		-- 008004: B240             MOV.W   #0x5a80,&WDTCTL_L
						   32773 => x"60",
						   32774 => x"80",		-- 008006: 805A            
						   32775 => x"5A",
						   32776 => x"CC",		-- 008008: CC01            
						   32777 => x"01",
						   32778 => x"34",		-- 00800a: 3440             MOV.W   #0x2000,R4
						   32779 => x"60",
						   32780 => x"00",		-- 00800c: 0020            
						   32781 => x"20",
						   32782 => x"05",		-- 00800e: 0544             MOV.W   R4,R5
						   32783 => x"64",
						   32784 => x"36",		-- 008010: 3640             MOV.W   #0x2004,R6
						   32785 => x"60",
						   32786 => x"04",		-- 008012: 0420            
						   32787 => x"20",
						   32788 => x"E2",		-- 008014: E2C3             BIC.B   #2,&P4DIR
						   32789 => x"E3",
						   32790 => x"25",		-- 008016: 2502            
						   32791 => x"02",
						   32792 => x"E2",		-- 008018: E2D3             BIS.B   #2,&P4REN
						   32793 => x"F3",
						   32794 => x"27",		-- 00801a: 2702            
						   32795 => x"02",
						   32796 => x"E2",		-- 00801c: E2D3             BIS.B   #2,&P4OUT
						   32797 => x"F3",
						   32798 => x"23",		-- 00801e: 2302            
						   32799 => x"02",
						   32800 => x"F2",		-- 008020: F2C3             BIC.B   #-1,&P4IFG
						   32801 => x"E3",
						   32802 => x"3D",		-- 008022: 3D02            
						   32803 => x"02",
						   32804 => x"E2",		-- 008024: E2D3             BIS.B   #2,&P4IES
						   32805 => x"F3",
						   32806 => x"39",		-- 008026: 3902            
						   32807 => x"02",
						   32808 => x"E2",		-- 008028: E2D3             BIS.B   #2,&P4IE
						   32809 => x"F3",
						   32810 => x"3B",		-- 00802a: 3B02            
						   32811 => x"02",
						   32812 => x"03",		-- 00802c: 0343             NOP     
						   32813 => x"63",
						   32814 => x"32",		-- 00802e: 32D2             EINT    
						   32815 => x"F2",
						   32816 => x"03",		-- 008030: 0343             NOP     
						   32817 => x"63",
						   32818 => x"32",		-- 008032: 32D2             EINT    
						   32819 => x"F2",
						   32820 => x"03",		-- 008034: 0343             NOP     
						   32821 => x"63",
						   32822 => x"32",		-- 008036: 32C2             DINT    
						   32823 => x"E2",
						   32824 => x"03",		-- 008038: 0343             NOP     
						   32825 => x"63",
						   32826 => x"D2",		-- 00803a: D2C3             BIC.B   #1,&PM5CTL0_L
						   32827 => x"E3",
						   32828 => x"30",		-- 00803c: 3001            
						   32829 => x"01",
						   32830 => x"17",		-- 00803e: 1742             MOV.W   &Con1,R7
						   32831 => x"62",
						   32832 => x"00",		-- 008040: 0020            
						   32833 => x"20",
						   32834 => x"18",		-- 008042: 1840             MOV.W   Con2,R8
						   32835 => x"60",
						   32836 => x"BE",		-- 008044: BE9F            
						   32837 => x"9F",
						   32838 => x"29",		-- 008046: 2944             MOV.W   @R4,R9
						   32839 => x"64",
						   32840 => x"3A",		-- 008048: 3A45             MOV.W   @R5+,R10
						   32841 => x"65",
						   32842 => x"3B",		-- 00804a: 3B45             MOV.W   @R5+,R11
						   32843 => x"65",
						   32844 => x"96",		-- 00804c: 9644             MOV.W   0x0002(R4),0x0004(R6)
						   32845 => x"64",
						   32846 => x"02",		-- 00804e: 0200            
						   32847 => x"00",
						   32848 => x"04",		-- 008050: 0400            
						   32849 => x"00",
						   32850 => x"34",		-- 008052: 3440             MOV.W   #0x2000,R4
						   32851 => x"60",
						   32852 => x"00",		-- 008054: 0020            
						   32853 => x"20",
						   32854 => x"80",		-- 008056: 8054             ADD.W   R4,Const2
						   32855 => x"74",
						   32856 => x"CA",		-- 008058: CA9F            
						   32857 => x"9F",
						   32858 => x"15",		-- 00805a: 1552             ADD.W   &Con1,R5
						   32859 => x"72",
						   32860 => x"00",		-- 00805c: 0020            
						   32861 => x"20",
						   32862 => x"34",		-- 00805e: 3440             MOV.W   #0x2000,R4
						   32863 => x"60",
						   32864 => x"00",		-- 008060: 0020            
						   32865 => x"20",
						   32866 => x"36",		-- 008062: 3640             MOV.W   #0x2004,R6
						   32867 => x"60",
						   32868 => x"04",		-- 008064: 0420            
						   32869 => x"20",
						   32870 => x"A6",		-- 008066: A654             ADD.W   @R4,0x0004(R6)
						   32871 => x"74",
						   32872 => x"04",		-- 008068: 0400            
						   32873 => x"00",
						   32874 => x"B0",		-- 00806a: B050             ADD.W   #0x2000,Var1
						   32875 => x"70",
						   32876 => x"00",		-- 00806c: 0020            
						   32877 => x"20",
						   32878 => x"96",		-- 00806e: 969F            
						   32879 => x"9F",
						   32880 => x"36",		-- 008070: 3655             ADD.W   @R5+,R6
						   32881 => x"75",
						   32882 => x"05",		-- 008072: 0564             ADDC.W  R4,R5
						   32883 => x"84",
						   32884 => x"80",		-- 008074: 8065             ADDC.W  R5,Const2
						   32885 => x"85",
						   32886 => x"AC",		-- 008076: AC9F            
						   32887 => x"9F",
						   32888 => x"15",		-- 008078: 1562             ADDC.W  &Con1,R5
						   32889 => x"82",
						   32890 => x"00",		-- 00807a: 0020            
						   32891 => x"20",
						   32892 => x"34",		-- 00807c: 3440             MOV.W   #0x2000,R4
						   32893 => x"60",
						   32894 => x"00",		-- 00807e: 0020            
						   32895 => x"20",
						   32896 => x"36",		-- 008080: 3640             MOV.W   #0x2004,R6
						   32897 => x"60",
						   32898 => x"04",		-- 008082: 0420            
						   32899 => x"20",
						   32900 => x"A6",		-- 008084: A664             ADDC.W  @R4,0x0004(R6)
						   32901 => x"84",
						   32902 => x"04",		-- 008086: 0400            
						   32903 => x"00",
						   32904 => x"B0",		-- 008088: B060             ADDC.W  #0x2000,Var1
						   32905 => x"80",
						   32906 => x"00",		-- 00808a: 0020            
						   32907 => x"20",
						   32908 => x"78",		-- 00808c: 789F            
						   32909 => x"9F",
						   32910 => x"36",		-- 00808e: 3665             ADDC.W  @R5+,R6
						   32911 => x"85",
						   32912 => x"12",		-- 008090: 12D3             SETC    
						   32913 => x"F3",
						   32914 => x"04",		-- 008092: 0463             ADC.W   R4
						   32915 => x"83",
						   32916 => x"80",		-- 008094: 8063             ADC.W   Const2
						   32917 => x"83",
						   32918 => x"8C",		-- 008096: 8C9F            
						   32919 => x"9F",
						   32920 => x"82",		-- 008098: 8263             ADC.W   &Con1
						   32921 => x"83",
						   32922 => x"00",		-- 00809a: 0020            
						   32923 => x"20",
						   32924 => x"B0",		-- 00809c: B040             MOV.W   #0x2000,Var1
						   32925 => x"60",
						   32926 => x"00",		-- 00809e: 0020            
						   32927 => x"20",
						   32928 => x"64",		-- 0080a0: 649F            
						   32929 => x"9F",
						   32930 => x"34",		-- 0080a2: 3440             MOV.W   #0x2000,R4
						   32931 => x"60",
						   32932 => x"00",		-- 0080a4: 0020            
						   32933 => x"20",
						   32934 => x"12",		-- 0080a6: 12D3             SETC    
						   32935 => x"F3",
						   32936 => x"80",		-- 0080a8: 8063             ADC.W   Var1
						   32937 => x"83",
						   32938 => x"5A",		-- 0080aa: 5A9F            
						   32939 => x"9F",
						   32940 => x"84",		-- 0080ac: 8463             ADC.W   0x0004(R4)
						   32941 => x"83",
						   32942 => x"04",		-- 0080ae: 0400            
						   32943 => x"00",
						   32944 => x"05",		-- 0080b0: 0584             SUB.W   R4,R5
						   32945 => x"A4",
						   32946 => x"80",		-- 0080b2: 8084             SUB.W   R4,Const2
						   32947 => x"A4",
						   32948 => x"6E",		-- 0080b4: 6E9F            
						   32949 => x"9F",
						   32950 => x"15",		-- 0080b6: 1582             SUB.W   &Con1,R5
						   32951 => x"A2",
						   32952 => x"00",		-- 0080b8: 0020            
						   32953 => x"20",
						   32954 => x"34",		-- 0080ba: 3440             MOV.W   #0x2000,R4
						   32955 => x"60",
						   32956 => x"00",		-- 0080bc: 0020            
						   32957 => x"20",
						   32958 => x"36",		-- 0080be: 3640             MOV.W   #0x2004,R6
						   32959 => x"60",
						   32960 => x"04",		-- 0080c0: 0420            
						   32961 => x"20",
						   32962 => x"A6",		-- 0080c2: A684             SUB.W   @R4,0x0004(R6)
						   32963 => x"A4",
						   32964 => x"04",		-- 0080c4: 0400            
						   32965 => x"00",
						   32966 => x"B0",		-- 0080c6: B080             SUB.W   #0x2000,Var1
						   32967 => x"A0",
						   32968 => x"00",		-- 0080c8: 0020            
						   32969 => x"20",
						   32970 => x"3A",		-- 0080ca: 3A9F            
						   32971 => x"9F",
						   32972 => x"36",		-- 0080cc: 3685             SUB.W   @R5+,R6
						   32973 => x"A5",
						   32974 => x"06",		-- 0080ce: 0675             SUBC.W  R5,R6
						   32975 => x"95",
						   32976 => x"80",		-- 0080d0: 8074             SUBC.W  R4,Const2
						   32977 => x"94",
						   32978 => x"50",		-- 0080d2: 509F            
						   32979 => x"9F",
						   32980 => x"15",		-- 0080d4: 1572             SUBC.W  &Con1,R5
						   32981 => x"92",
						   32982 => x"00",		-- 0080d6: 0020            
						   32983 => x"20",
						   32984 => x"34",		-- 0080d8: 3440             MOV.W   #0x2000,R4
						   32985 => x"60",
						   32986 => x"00",		-- 0080da: 0020            
						   32987 => x"20",
						   32988 => x"36",		-- 0080dc: 3640             MOV.W   #0x2004,R6
						   32989 => x"60",
						   32990 => x"04",		-- 0080de: 0420            
						   32991 => x"20",
						   32992 => x"A6",		-- 0080e0: A674             SUBC.W  @R4,0x0004(R6)
						   32993 => x"94",
						   32994 => x"04",		-- 0080e2: 0400            
						   32995 => x"00",
						   32996 => x"B0",		-- 0080e4: B070             SUBC.W  #0x2000,Var1
						   32997 => x"90",
						   32998 => x"00",		-- 0080e6: 0020            
						   32999 => x"20",
						   33000 => x"1C",		-- 0080e8: 1C9F            
						   33001 => x"9F",
						   33002 => x"36",		-- 0080ea: 3675             SUBC.W  @R5+,R6
						   33003 => x"95",
						   33004 => x"12",		-- 0080ec: 12D3             SETC    
						   33005 => x"F3",
						   33006 => x"04",		-- 0080ee: 0473             SBC.W   R4
						   33007 => x"93",
						   33008 => x"80",		-- 0080f0: 8073             SBC.W   Const2
						   33009 => x"93",
						   33010 => x"30",		-- 0080f2: 309F            
						   33011 => x"9F",
						   33012 => x"82",		-- 0080f4: 8273             SBC.W   &Con1
						   33013 => x"93",
						   33014 => x"00",		-- 0080f6: 0020            
						   33015 => x"20",
						   33016 => x"B0",		-- 0080f8: B040             MOV.W   #0x2000,Var1
						   33017 => x"60",
						   33018 => x"00",		-- 0080fa: 0020            
						   33019 => x"20",
						   33020 => x"08",		-- 0080fc: 089F            
						   33021 => x"9F",
						   33022 => x"34",		-- 0080fe: 3440             MOV.W   #0x2000,R4
						   33023 => x"60",
						   33024 => x"00",		-- 008100: 0020            
						   33025 => x"20",
						   33026 => x"12",		-- 008102: 12D3             SETC    
						   33027 => x"F3",
						   33028 => x"80",		-- 008104: 8073             SBC.W   Var1
						   33029 => x"93",
						   33030 => x"FE",		-- 008106: FE9E            
						   33031 => x"9E",
						   33032 => x"84",		-- 008108: 8473             SBC.W   0x0004(R4)
						   33033 => x"93",
						   33034 => x"04",		-- 00810a: 0400            
						   33035 => x"00",
						   33036 => x"12",		-- 00810c: 12D3             SETC    
						   33037 => x"F3",
						   33038 => x"05",		-- 00810e: 05A4             DADD.W  R4,R5
						   33039 => x"C4",
						   33040 => x"80",		-- 008110: 80A4             DADD.W  R4,Const2
						   33041 => x"C4",
						   33042 => x"10",		-- 008112: 109F            
						   33043 => x"9F",
						   33044 => x"15",		-- 008114: 15A2             DADD.W  &Con1,R5
						   33045 => x"C2",
						   33046 => x"00",		-- 008116: 0020            
						   33047 => x"20",
						   33048 => x"34",		-- 008118: 3440             MOV.W   #0x2000,R4
						   33049 => x"60",
						   33050 => x"00",		-- 00811a: 0020            
						   33051 => x"20",
						   33052 => x"36",		-- 00811c: 3640             MOV.W   #0x2004,R6
						   33053 => x"60",
						   33054 => x"04",		-- 00811e: 0420            
						   33055 => x"20",
						   33056 => x"12",		-- 008120: 12D3             SETC    
						   33057 => x"F3",
						   33058 => x"A6",		-- 008122: A6A4             DADD.W  @R4,0x0004(R6)
						   33059 => x"C4",
						   33060 => x"04",		-- 008124: 0400            
						   33061 => x"00",
						   33062 => x"B0",		-- 008126: B0A0             DADD.W  #0x2000,Var1
						   33063 => x"C0",
						   33064 => x"00",		-- 008128: 0020            
						   33065 => x"20",
						   33066 => x"DA",		-- 00812a: DA9E            
						   33067 => x"9E",
						   33068 => x"36",		-- 00812c: 36A5             DADD.W  @R5+,R6
						   33069 => x"C5",
						   33070 => x"12",		-- 00812e: 12D3             SETC    
						   33071 => x"F3",
						   33072 => x"04",		-- 008130: 04A3             DADC.W  R4
						   33073 => x"C3",
						   33074 => x"80",		-- 008132: 80A3             DADC.W  Const2
						   33075 => x"C3",
						   33076 => x"EE",		-- 008134: EE9E            
						   33077 => x"9E",
						   33078 => x"82",		-- 008136: 82A3             DADC.W  &Con1
						   33079 => x"C3",
						   33080 => x"00",		-- 008138: 0020            
						   33081 => x"20",
						   33082 => x"B0",		-- 00813a: B040             MOV.W   #0x2000,Var1
						   33083 => x"60",
						   33084 => x"00",		-- 00813c: 0020            
						   33085 => x"20",
						   33086 => x"C6",		-- 00813e: C69E            
						   33087 => x"9E",
						   33088 => x"34",		-- 008140: 3440             MOV.W   #0x2000,R4
						   33089 => x"60",
						   33090 => x"00",		-- 008142: 0020            
						   33091 => x"20",
						   33092 => x"12",		-- 008144: 12D3             SETC    
						   33093 => x"F3",
						   33094 => x"80",		-- 008146: 80A3             DADC.W  Var1
						   33095 => x"C3",
						   33096 => x"BC",		-- 008148: BC9E            
						   33097 => x"9E",
						   33098 => x"84",		-- 00814a: 84A3             DADC.W  0x0004(R4)
						   33099 => x"C3",
						   33100 => x"04",		-- 00814c: 0400            
						   33101 => x"00",
						   33102 => x"14",		-- 00814e: 1453             INC.W   R4
						   33103 => x"73",
						   33104 => x"90",		-- 008150: 9053             INC.W   Const2
						   33105 => x"73",
						   33106 => x"D0",		-- 008152: D09E            
						   33107 => x"9E",
						   33108 => x"92",		-- 008154: 9253             INC.W   &Con1
						   33109 => x"73",
						   33110 => x"00",		-- 008156: 0020            
						   33111 => x"20",
						   33112 => x"B0",		-- 008158: B040             MOV.W   #0x2000,Var1
						   33113 => x"60",
						   33114 => x"00",		-- 00815a: 0020            
						   33115 => x"20",
						   33116 => x"A8",		-- 00815c: A89E            
						   33117 => x"9E",
						   33118 => x"34",		-- 00815e: 3440             MOV.W   #0x2000,R4
						   33119 => x"60",
						   33120 => x"00",		-- 008160: 0020            
						   33121 => x"20",
						   33122 => x"90",		-- 008162: 9053             INC.W   Var1
						   33123 => x"73",
						   33124 => x"A0",		-- 008164: A09E            
						   33125 => x"9E",
						   33126 => x"94",		-- 008166: 9453             INC.W   0x0004(R4)
						   33127 => x"73",
						   33128 => x"04",		-- 008168: 0400            
						   33129 => x"00",
						   33130 => x"24",		-- 00816a: 2453             INCD.W  R4
						   33131 => x"73",
						   33132 => x"A0",		-- 00816c: A053             INCD.W  Const2
						   33133 => x"73",
						   33134 => x"B4",		-- 00816e: B49E            
						   33135 => x"9E",
						   33136 => x"A2",		-- 008170: A253             INCD.W  &Con1
						   33137 => x"73",
						   33138 => x"00",		-- 008172: 0020            
						   33139 => x"20",
						   33140 => x"B0",		-- 008174: B040             MOV.W   #0x2000,Var1
						   33141 => x"60",
						   33142 => x"00",		-- 008176: 0020            
						   33143 => x"20",
						   33144 => x"8C",		-- 008178: 8C9E            
						   33145 => x"9E",
						   33146 => x"34",		-- 00817a: 3440             MOV.W   #0x2000,R4
						   33147 => x"60",
						   33148 => x"00",		-- 00817c: 0020            
						   33149 => x"20",
						   33150 => x"A0",		-- 00817e: A053             INCD.W  Var1
						   33151 => x"73",
						   33152 => x"84",		-- 008180: 849E            
						   33153 => x"9E",
						   33154 => x"A4",		-- 008182: A453             INCD.W  0x0004(R4)
						   33155 => x"73",
						   33156 => x"04",		-- 008184: 0400            
						   33157 => x"00",
						   33158 => x"14",		-- 008186: 1483             DEC.W   R4
						   33159 => x"A3",
						   33160 => x"90",		-- 008188: 9083             DEC.W   Const2
						   33161 => x"A3",
						   33162 => x"98",		-- 00818a: 989E            
						   33163 => x"9E",
						   33164 => x"92",		-- 00818c: 9283             DEC.W   &Con1
						   33165 => x"A3",
						   33166 => x"00",		-- 00818e: 0020            
						   33167 => x"20",
						   33168 => x"B0",		-- 008190: B040             MOV.W   #0x2000,Var1
						   33169 => x"60",
						   33170 => x"00",		-- 008192: 0020            
						   33171 => x"20",
						   33172 => x"70",		-- 008194: 709E            
						   33173 => x"9E",
						   33174 => x"34",		-- 008196: 3440             MOV.W   #0x2000,R4
						   33175 => x"60",
						   33176 => x"00",		-- 008198: 0020            
						   33177 => x"20",
						   33178 => x"90",		-- 00819a: 9083             DEC.W   Var1
						   33179 => x"A3",
						   33180 => x"68",		-- 00819c: 689E            
						   33181 => x"9E",
						   33182 => x"94",		-- 00819e: 9483             DEC.W   0x0004(R4)
						   33183 => x"A3",
						   33184 => x"04",		-- 0081a0: 0400            
						   33185 => x"00",
						   33186 => x"24",		-- 0081a2: 2483             DECD.W  R4
						   33187 => x"A3",
						   33188 => x"A0",		-- 0081a4: A083             DECD.W  Const2
						   33189 => x"A3",
						   33190 => x"7C",		-- 0081a6: 7C9E            
						   33191 => x"9E",
						   33192 => x"A2",		-- 0081a8: A283             DECD.W  &Con1
						   33193 => x"A3",
						   33194 => x"00",		-- 0081aa: 0020            
						   33195 => x"20",
						   33196 => x"B0",		-- 0081ac: B040             MOV.W   #0x2000,Var1
						   33197 => x"60",
						   33198 => x"00",		-- 0081ae: 0020            
						   33199 => x"20",
						   33200 => x"54",		-- 0081b0: 549E            
						   33201 => x"9E",
						   33202 => x"34",		-- 0081b2: 3440             MOV.W   #0x2000,R4
						   33203 => x"60",
						   33204 => x"00",		-- 0081b4: 0020            
						   33205 => x"20",
						   33206 => x"A0",		-- 0081b6: A083             DECD.W  Var1
						   33207 => x"A3",
						   33208 => x"4C",		-- 0081b8: 4C9E            
						   33209 => x"9E",
						   33210 => x"A4",		-- 0081ba: A483             DECD.W  0x0004(R4)
						   33211 => x"A3",
						   33212 => x"04",		-- 0081bc: 0400            
						   33213 => x"00",
						   33214 => x"74",		-- 0081be: 7440             MOV.B   #0x004e,R4
						   33215 => x"60",
						   33216 => x"4E",		-- 0081c0: 4E00            
						   33217 => x"00",
						   33218 => x"74",		-- 0081c2: 74E3             INV.B   R4
						   33219 => x"03",
						   33220 => x"34",		-- 0081c4: 3440             MOV.W   #0x2032,R4
						   33221 => x"60",
						   33222 => x"32",		-- 0081c6: 3220            
						   33223 => x"20",
						   33224 => x"34",		-- 0081c8: 34E3             INV.W   R4
						   33225 => x"03",
						   33226 => x"B2",		-- 0081ca: B2E3             INV.W   &Const1
						   33227 => x"03",
						   33228 => x"20",		-- 0081cc: 2020            
						   33229 => x"20",
						   33230 => x"B0",		-- 0081ce: B0E3             INV.W   Const10
						   33231 => x"03",
						   33232 => x"62",		-- 0081d0: 629E            
						   33233 => x"9E",
						   33234 => x"34",		-- 0081d2: 3440             MOV.W   #0x2032,R4
						   33235 => x"60",
						   33236 => x"32",		-- 0081d4: 3220            
						   33237 => x"20",
						   33238 => x"B4",		-- 0081d6: B4E3             INV.W   0x0002(R4)
						   33239 => x"03",
						   33240 => x"02",		-- 0081d8: 0200            
						   33241 => x"00",
						   33242 => x"74",		-- 0081da: 7440             MOV.B   #0x00aa,R4
						   33243 => x"60",
						   33244 => x"AA",		-- 0081dc: AA00            
						   33245 => x"00",
						   33246 => x"74",		-- 0081de: 74F0             AND.B   #0x000f,R4
						   33247 => x"10",
						   33248 => x"0F",		-- 0081e0: 0F00            
						   33249 => x"00",
						   33250 => x"05",		-- 0081e2: 05F4             AND.W   R4,R5
						   33251 => x"14",
						   33252 => x"80",		-- 0081e4: 80F4             AND.W   R4,Const2
						   33253 => x"14",
						   33254 => x"3C",		-- 0081e6: 3C9E            
						   33255 => x"9E",
						   33256 => x"15",		-- 0081e8: 15F2             AND.W   &Con1,R5
						   33257 => x"12",
						   33258 => x"00",		-- 0081ea: 0020            
						   33259 => x"20",
						   33260 => x"34",		-- 0081ec: 3440             MOV.W   #0x2000,R4
						   33261 => x"60",
						   33262 => x"00",		-- 0081ee: 0020            
						   33263 => x"20",
						   33264 => x"36",		-- 0081f0: 3640             MOV.W   #0x2004,R6
						   33265 => x"60",
						   33266 => x"04",		-- 0081f2: 0420            
						   33267 => x"20",
						   33268 => x"A6",		-- 0081f4: A6F4             AND.W   @R4,0x0004(R6)
						   33269 => x"14",
						   33270 => x"04",		-- 0081f6: 0400            
						   33271 => x"00",
						   33272 => x"B0",		-- 0081f8: B0F0             AND.W   #0x2000,Var1
						   33273 => x"10",
						   33274 => x"00",		-- 0081fa: 0020            
						   33275 => x"20",
						   33276 => x"08",		-- 0081fc: 089E            
						   33277 => x"9E",
						   33278 => x"36",		-- 0081fe: 36F5             AND.W   @R5+,R6
						   33279 => x"15",
						   33280 => x"74",		-- 008200: 7440             MOV.B   #0x00aa,R4
						   33281 => x"60",
						   33282 => x"AA",		-- 008202: AA00            
						   33283 => x"00",
						   33284 => x"74",		-- 008204: 74D0             BIS.B   #0x0249,R4
						   33285 => x"F0",
						   33286 => x"49",		-- 008206: 4902            
						   33287 => x"02",
						   33288 => x"05",		-- 008208: 05D4             BIS.W   R4,R5
						   33289 => x"F4",
						   33290 => x"80",		-- 00820a: 80D4             BIS.W   R4,Const2
						   33291 => x"F4",
						   33292 => x"16",		-- 00820c: 169E            
						   33293 => x"9E",
						   33294 => x"15",		-- 00820e: 15D2             BIS.W   &Con1,R5
						   33295 => x"F2",
						   33296 => x"00",		-- 008210: 0020            
						   33297 => x"20",
						   33298 => x"34",		-- 008212: 34D0             BIS.W   #0x2000,R4
						   33299 => x"F0",
						   33300 => x"00",		-- 008214: 0020            
						   33301 => x"20",
						   33302 => x"36",		-- 008216: 36D0             BIS.W   #0x2004,R6
						   33303 => x"F0",
						   33304 => x"04",		-- 008218: 0420            
						   33305 => x"20",
						   33306 => x"A6",		-- 00821a: A6D4             BIS.W   @R4,0x0004(R6)
						   33307 => x"F4",
						   33308 => x"04",		-- 00821c: 0400            
						   33309 => x"00",
						   33310 => x"B0",		-- 00821e: B0D0             BIS.W   #0x2000,Var1
						   33311 => x"F0",
						   33312 => x"00",		-- 008220: 0020            
						   33313 => x"20",
						   33314 => x"E2",		-- 008222: E29D            
						   33315 => x"9D",
						   33316 => x"36",		-- 008224: 36D5             BIS.W   @R5+,R6
						   33317 => x"F5",
						   33318 => x"74",		-- 008226: 7440             MOV.B   #0x00aa,R4
						   33319 => x"60",
						   33320 => x"AA",		-- 008228: AA00            
						   33321 => x"00",
						   33322 => x"74",		-- 00822a: 74E0             XOR.B   #0x0055,R4
						   33323 => x"00",
						   33324 => x"55",		-- 00822c: 5500            
						   33325 => x"00",
						   33326 => x"06",		-- 00822e: 06E5             XOR.W   R5,R6
						   33327 => x"05",
						   33328 => x"80",		-- 008230: 80E4             XOR.W   R4,Const2
						   33329 => x"04",
						   33330 => x"F0",		-- 008232: F09D            
						   33331 => x"9D",
						   33332 => x"15",		-- 008234: 15E2             XOR.W   &Con1,R5
						   33333 => x"02",
						   33334 => x"00",		-- 008236: 0020            
						   33335 => x"20",
						   33336 => x"34",		-- 008238: 3440             MOV.W   #0x2000,R4
						   33337 => x"60",
						   33338 => x"00",		-- 00823a: 0020            
						   33339 => x"20",
						   33340 => x"36",		-- 00823c: 3640             MOV.W   #0x2004,R6
						   33341 => x"60",
						   33342 => x"04",		-- 00823e: 0420            
						   33343 => x"20",
						   33344 => x"A6",		-- 008240: A6E4             XOR.W   @R4,0x0004(R6)
						   33345 => x"04",
						   33346 => x"04",		-- 008242: 0400            
						   33347 => x"00",
						   33348 => x"B0",		-- 008244: B0E0             XOR.W   #0x2000,Var1
						   33349 => x"00",
						   33350 => x"00",		-- 008246: 0020            
						   33351 => x"20",
						   33352 => x"BC",		-- 008248: BC9D            
						   33353 => x"9D",
						   33354 => x"36",		-- 00824a: 36E5             XOR.W   @R5+,R6
						   33355 => x"05",
						   33356 => x"74",		-- 00824c: 7440             MOV.B   #0x00aa,R4
						   33357 => x"60",
						   33358 => x"AA",		-- 00824e: AA00            
						   33359 => x"00",
						   33360 => x"74",		-- 008250: 74D0             BIS.B   #0x0249,R4
						   33361 => x"F0",
						   33362 => x"49",		-- 008252: 4902            
						   33363 => x"02",
						   33364 => x"05",		-- 008254: 05D4             BIS.W   R4,R5
						   33365 => x"F4",
						   33366 => x"80",		-- 008256: 80D4             BIS.W   R4,Const2
						   33367 => x"F4",
						   33368 => x"CA",		-- 008258: CA9D            
						   33369 => x"9D",
						   33370 => x"15",		-- 00825a: 15D2             BIS.W   &Con1,R5
						   33371 => x"F2",
						   33372 => x"00",		-- 00825c: 0020            
						   33373 => x"20",
						   33374 => x"34",		-- 00825e: 3440             MOV.W   #0x2000,R4
						   33375 => x"60",
						   33376 => x"00",		-- 008260: 0020            
						   33377 => x"20",
						   33378 => x"36",		-- 008262: 3640             MOV.W   #0x2004,R6
						   33379 => x"60",
						   33380 => x"04",		-- 008264: 0420            
						   33381 => x"20",
						   33382 => x"A6",		-- 008266: A6D4             BIS.W   @R4,0x0004(R6)
						   33383 => x"F4",
						   33384 => x"04",		-- 008268: 0400            
						   33385 => x"00",
						   33386 => x"B0",		-- 00826a: B0D0             BIS.W   #0x2000,Var1
						   33387 => x"F0",
						   33388 => x"00",		-- 00826c: 0020            
						   33389 => x"20",
						   33390 => x"96",		-- 00826e: 969D            
						   33391 => x"9D",
						   33392 => x"36",		-- 008270: 36D5             BIS.W   @R5+,R6
						   33393 => x"F5",
						   33394 => x"74",		-- 008272: 7440             MOV.B   #0x00aa,R4
						   33395 => x"60",
						   33396 => x"AA",		-- 008274: AA00            
						   33397 => x"00",
						   33398 => x"74",		-- 008276: 74C0             BIC.B   #0x0018,R4
						   33399 => x"E0",
						   33400 => x"18",		-- 008278: 1800            
						   33401 => x"00",
						   33402 => x"05",		-- 00827a: 05C4             BIC.W   R4,R5
						   33403 => x"E4",
						   33404 => x"80",		-- 00827c: 80C4             BIC.W   R4,Const2
						   33405 => x"E4",
						   33406 => x"A4",		-- 00827e: A49D            
						   33407 => x"9D",
						   33408 => x"15",		-- 008280: 15C2             BIC.W   &Con1,R5
						   33409 => x"E2",
						   33410 => x"00",		-- 008282: 0020            
						   33411 => x"20",
						   33412 => x"34",		-- 008284: 3440             MOV.W   #0x2000,R4
						   33413 => x"60",
						   33414 => x"00",		-- 008286: 0020            
						   33415 => x"20",
						   33416 => x"36",		-- 008288: 3640             MOV.W   #0x2004,R6
						   33417 => x"60",
						   33418 => x"04",		-- 00828a: 0420            
						   33419 => x"20",
						   33420 => x"A6",		-- 00828c: A6C4             BIC.W   @R4,0x0004(R6)
						   33421 => x"E4",
						   33422 => x"04",		-- 00828e: 0400            
						   33423 => x"00",
						   33424 => x"B0",		-- 008290: B0C0             BIC.W   #0x2000,Var1
						   33425 => x"E0",
						   33426 => x"00",		-- 008292: 0020            
						   33427 => x"20",
						   33428 => x"70",		-- 008294: 709D            
						   33429 => x"9D",
						   33430 => x"36",		-- 008296: 36C5             BIC.W   @R5+,R6
						   33431 => x"E5",
						   33432 => x"74",		-- 008298: 7440             MOV.B   #0x00aa,R4
						   33433 => x"60",
						   33434 => x"AA",		-- 00829a: AA00            
						   33435 => x"00",
						   33436 => x"74",		-- 00829c: 74B0             BIT.B   #0x0018,R4
						   33437 => x"D0",
						   33438 => x"18",		-- 00829e: 1800            
						   33439 => x"00",
						   33440 => x"05",		-- 0082a0: 05B4             BIT.W   R4,R5
						   33441 => x"D4",
						   33442 => x"80",		-- 0082a2: 80B4             BIT.W   R4,Const2
						   33443 => x"D4",
						   33444 => x"7E",		-- 0082a4: 7E9D            
						   33445 => x"9D",
						   33446 => x"15",		-- 0082a6: 15B2             BIT.W   &Con1,R5
						   33447 => x"D2",
						   33448 => x"00",		-- 0082a8: 0020            
						   33449 => x"20",
						   33450 => x"34",		-- 0082aa: 3440             MOV.W   #0x2000,R4
						   33451 => x"60",
						   33452 => x"00",		-- 0082ac: 0020            
						   33453 => x"20",
						   33454 => x"36",		-- 0082ae: 3640             MOV.W   #0x2004,R6
						   33455 => x"60",
						   33456 => x"04",		-- 0082b0: 0420            
						   33457 => x"20",
						   33458 => x"A6",		-- 0082b2: A6B4             BIT.W   @R4,0x0004(R6)
						   33459 => x"D4",
						   33460 => x"04",		-- 0082b4: 0400            
						   33461 => x"00",
						   33462 => x"B0",		-- 0082b6: B0B0             BIT.W   #0x2000,Var1
						   33463 => x"D0",
						   33464 => x"00",		-- 0082b8: 0020            
						   33465 => x"20",
						   33466 => x"4A",		-- 0082ba: 4A9D            
						   33467 => x"9D",
						   33468 => x"36",		-- 0082bc: 36B5             BIT.W   @R5+,R6
						   33469 => x"D5",
						   33470 => x"75",		-- 0082be: 7540             MOV.B   #0x0063,R5
						   33471 => x"60",
						   33472 => x"63",		-- 0082c0: 6300            
						   33473 => x"00",
						   33474 => x"75",		-- 0082c2: 7590             CMP.B   #0x0063,R5
						   33475 => x"B0",
						   33476 => x"63",		-- 0082c4: 6300            
						   33477 => x"00",
						   33478 => x"75",		-- 0082c6: 7590             CMP.B   #0x004d,R5
						   33479 => x"B0",
						   33480 => x"4D",		-- 0082c8: 4D00            
						   33481 => x"00",
						   33482 => x"05",		-- 0082ca: 0594             CMP.W   R4,R5
						   33483 => x"B4",
						   33484 => x"80",		-- 0082cc: 8094             CMP.W   R4,Const2
						   33485 => x"B4",
						   33486 => x"54",		-- 0082ce: 549D            
						   33487 => x"9D",
						   33488 => x"15",		-- 0082d0: 1592             CMP.W   &Con1,R5
						   33489 => x"B2",
						   33490 => x"00",		-- 0082d2: 0020            
						   33491 => x"20",
						   33492 => x"34",		-- 0082d4: 3440             MOV.W   #0x2000,R4
						   33493 => x"60",
						   33494 => x"00",		-- 0082d6: 0020            
						   33495 => x"20",
						   33496 => x"36",		-- 0082d8: 3640             MOV.W   #0x2004,R6
						   33497 => x"60",
						   33498 => x"04",		-- 0082da: 0420            
						   33499 => x"20",
						   33500 => x"A6",		-- 0082dc: A694             CMP.W   @R4,0x0004(R6)
						   33501 => x"B4",
						   33502 => x"04",		-- 0082de: 0400            
						   33503 => x"00",
						   33504 => x"B0",		-- 0082e0: B090             CMP.W   #0x2000,Var1
						   33505 => x"B0",
						   33506 => x"00",		-- 0082e2: 0020            
						   33507 => x"20",
						   33508 => x"20",		-- 0082e4: 209D            
						   33509 => x"9D",
						   33510 => x"36",		-- 0082e6: 3695             CMP.W   @R5+,R6
						   33511 => x"B5",
						   33512 => x"77",		-- 0082e8: 7740             MOV.B   #0xff9d,R7
						   33513 => x"60",
						   33514 => x"9D",		-- 0082ea: 9DFF            
						   33515 => x"FF",
						   33516 => x"46",		-- 0082ec: 4643             CLR.B   R6
						   33517 => x"63",
						   33518 => x"46",		-- 0082ee: 4693             TST.B   R6
						   33519 => x"B3",
						   33520 => x"47",		-- 0082f0: 4793             TST.B   R7
						   33521 => x"B3",
						   33522 => x"04",		-- 0082f2: 0493             TST.W   R4
						   33523 => x"B3",
						   33524 => x"80",		-- 0082f4: 8093             TST.W   Const2
						   33525 => x"B3",
						   33526 => x"2C",		-- 0082f6: 2C9D            
						   33527 => x"9D",
						   33528 => x"82",		-- 0082f8: 8293             TST.W   &Con1
						   33529 => x"B3",
						   33530 => x"00",		-- 0082fa: 0020            
						   33531 => x"20",
						   33532 => x"B0",		-- 0082fc: B040             MOV.W   #0x2000,Var1
						   33533 => x"60",
						   33534 => x"00",		-- 0082fe: 0020            
						   33535 => x"20",
						   33536 => x"04",		-- 008300: 049D            
						   33537 => x"9D",
						   33538 => x"34",		-- 008302: 3440             MOV.W   #0x2000,R4
						   33539 => x"60",
						   33540 => x"00",		-- 008304: 0020            
						   33541 => x"20",
						   33542 => x"80",		-- 008306: 8093             TST.W   Var1
						   33543 => x"B3",
						   33544 => x"FC",		-- 008308: FC9C            
						   33545 => x"9C",
						   33546 => x"84",		-- 00830a: 8493             TST.W   0x0004(R4)
						   33547 => x"B3",
						   33548 => x"04",		-- 00830c: 0400            
						   33549 => x"00",
						   33550 => x"54",		-- 00830e: 5443             MOV.B   #1,R4
						   33551 => x"63",
						   33552 => x"44",		-- 008310: 4454             RLA.B   R4
						   33553 => x"74",
						   33554 => x"44",		-- 008312: 4454             RLA.B   R4
						   33555 => x"74",
						   33556 => x"04",		-- 008314: 0454             RLA.W   R4
						   33557 => x"74",
						   33558 => x"90",		-- 008316: 9050             ADD.W   Const2,Const2
						   33559 => x"70",
						   33560 => x"0A",		-- 008318: 0A9D            
						   33561 => x"9D",
						   33562 => x"08",		-- 00831a: 089D            
						   33563 => x"9D",
						   33564 => x"92",		-- 00831c: 9252             RLA.W   &Con1
						   33565 => x"72",
						   33566 => x"00",		-- 00831e: 0020            
						   33567 => x"20",
						   33568 => x"00",		-- 008320: 0020            
						   33569 => x"20",
						   33570 => x"B0",		-- 008322: B040             MOV.W   #0x2000,Var1
						   33571 => x"60",
						   33572 => x"00",		-- 008324: 0020            
						   33573 => x"20",
						   33574 => x"DE",		-- 008326: DE9C            
						   33575 => x"9C",
						   33576 => x"34",		-- 008328: 3440             MOV.W   #0x2000,R4
						   33577 => x"60",
						   33578 => x"00",		-- 00832a: 0020            
						   33579 => x"20",
						   33580 => x"90",		-- 00832c: 9050             ADD.W   Var1,Var1
						   33581 => x"70",
						   33582 => x"D6",		-- 00832e: D69C            
						   33583 => x"9C",
						   33584 => x"D4",		-- 008330: D49C            
						   33585 => x"9C",
						   33586 => x"94",		-- 008332: 9454             RLA.W   0x0004(R4)
						   33587 => x"74",
						   33588 => x"04",		-- 008334: 0400            
						   33589 => x"00",
						   33590 => x"04",		-- 008336: 0400            
						   33591 => x"00",
						   33592 => x"74",		-- 008338: 7440             MOV.B   #0x0020,R4
						   33593 => x"60",
						   33594 => x"20",		-- 00833a: 2000            
						   33595 => x"00",
						   33596 => x"44",		-- 00833c: 4411             RRA.B   R4
						   33597 => x"31",
						   33598 => x"44",		-- 00833e: 4411             RRA.B   R4
						   33599 => x"31",
						   33600 => x"04",		-- 008340: 0411             RRA     R4
						   33601 => x"31",
						   33602 => x"10",		-- 008342: 1011             RRA     Const2
						   33603 => x"31",
						   33604 => x"DE",		-- 008344: DE9C            
						   33605 => x"9C",
						   33606 => x"12",		-- 008346: 1211             RRA     &Con1
						   33607 => x"31",
						   33608 => x"00",		-- 008348: 0020            
						   33609 => x"20",
						   33610 => x"B0",		-- 00834a: B040             MOV.W   #0x2000,Var1
						   33611 => x"60",
						   33612 => x"00",		-- 00834c: 0020            
						   33613 => x"20",
						   33614 => x"B6",		-- 00834e: B69C            
						   33615 => x"9C",
						   33616 => x"34",		-- 008350: 3440             MOV.W   #0x2000,R4
						   33617 => x"60",
						   33618 => x"00",		-- 008352: 0020            
						   33619 => x"20",
						   33620 => x"10",		-- 008354: 1011             RRA     Var1
						   33621 => x"31",
						   33622 => x"AE",		-- 008356: AE9C            
						   33623 => x"9C",
						   33624 => x"14",		-- 008358: 1411             RRA     0x0004(R4)
						   33625 => x"31",
						   33626 => x"04",		-- 00835a: 0400            
						   33627 => x"00",
						   33628 => x"12",		-- 00835c: 12C3             CLRC    
						   33629 => x"E3",
						   33630 => x"77",		-- 00835e: 7740             MOV.B   #0x0080,R7
						   33631 => x"60",
						   33632 => x"80",		-- 008360: 8000            
						   33633 => x"00",
						   33634 => x"47",		-- 008362: 4767             RLC.B   R7
						   33635 => x"87",
						   33636 => x"47",		-- 008364: 4767             RLC.B   R7
						   33637 => x"87",
						   33638 => x"04",		-- 008366: 0464             RLC.W   R4
						   33639 => x"84",
						   33640 => x"90",		-- 008368: 9060             ADDC.W  Const2,Const2
						   33641 => x"80",
						   33642 => x"B8",		-- 00836a: B89C            
						   33643 => x"9C",
						   33644 => x"B6",		-- 00836c: B69C            
						   33645 => x"9C",
						   33646 => x"92",		-- 00836e: 9262             RLC.W   &Con1
						   33647 => x"82",
						   33648 => x"00",		-- 008370: 0020            
						   33649 => x"20",
						   33650 => x"00",		-- 008372: 0020            
						   33651 => x"20",
						   33652 => x"B0",		-- 008374: B040             MOV.W   #0x2000,Var1
						   33653 => x"60",
						   33654 => x"00",		-- 008376: 0020            
						   33655 => x"20",
						   33656 => x"8C",		-- 008378: 8C9C            
						   33657 => x"9C",
						   33658 => x"34",		-- 00837a: 3440             MOV.W   #0x2000,R4
						   33659 => x"60",
						   33660 => x"00",		-- 00837c: 0020            
						   33661 => x"20",
						   33662 => x"90",		-- 00837e: 9060             ADDC.W  Var1,Var1
						   33663 => x"80",
						   33664 => x"84",		-- 008380: 849C            
						   33665 => x"9C",
						   33666 => x"82",		-- 008382: 829C            
						   33667 => x"9C",
						   33668 => x"94",		-- 008384: 9464             RLC.W   0x0004(R4)
						   33669 => x"84",
						   33670 => x"04",		-- 008386: 0400            
						   33671 => x"00",
						   33672 => x"04",		-- 008388: 0400            
						   33673 => x"00",
						   33674 => x"12",		-- 00838a: 12C3             CLRC    
						   33675 => x"E3",
						   33676 => x"58",		-- 00838c: 5843             MOV.B   #1,R8
						   33677 => x"63",
						   33678 => x"48",		-- 00838e: 4810             RRC.B   R8
						   33679 => x"30",
						   33680 => x"48",		-- 008390: 4810             RRC.B   R8
						   33681 => x"30",
						   33682 => x"04",		-- 008392: 0410             RRC     R4
						   33683 => x"30",
						   33684 => x"10",		-- 008394: 1010             RRC     Const2
						   33685 => x"30",
						   33686 => x"8C",		-- 008396: 8C9C            
						   33687 => x"9C",
						   33688 => x"12",		-- 008398: 1210             RRC     &Con1
						   33689 => x"30",
						   33690 => x"00",		-- 00839a: 0020            
						   33691 => x"20",
						   33692 => x"B0",		-- 00839c: B040             MOV.W   #0x2000,Var1
						   33693 => x"60",
						   33694 => x"00",		-- 00839e: 0020            
						   33695 => x"20",
						   33696 => x"64",		-- 0083a0: 649C            
						   33697 => x"9C",
						   33698 => x"34",		-- 0083a2: 3440             MOV.W   #0x2000,R4
						   33699 => x"60",
						   33700 => x"00",		-- 0083a4: 0020            
						   33701 => x"20",
						   33702 => x"10",		-- 0083a6: 1010             RRC     Var1
						   33703 => x"30",
						   33704 => x"5C",		-- 0083a8: 5C9C            
						   33705 => x"9C",
						   33706 => x"14",		-- 0083aa: 1410             RRC     0x0004(R4)
						   33707 => x"30",
						   33708 => x"04",		-- 0083ac: 0400            
						   33709 => x"00",
						   33710 => x"34",		-- 0083ae: 3440             MOV.W   #0x00ff,R4
						   33711 => x"60",
						   33712 => x"FF",		-- 0083b0: FF00            
						   33713 => x"00",
						   33714 => x"84",		-- 0083b2: 8410             SWPB    R4
						   33715 => x"30",
						   33716 => x"90",		-- 0083b4: 9010             SWPB    Const2
						   33717 => x"30",
						   33718 => x"6C",		-- 0083b6: 6C9C            
						   33719 => x"9C",
						   33720 => x"92",		-- 0083b8: 9210             SWPB    &Con1
						   33721 => x"30",
						   33722 => x"00",		-- 0083ba: 0020            
						   33723 => x"20",
						   33724 => x"B0",		-- 0083bc: B040             MOV.W   #0x2000,Var1
						   33725 => x"60",
						   33726 => x"00",		-- 0083be: 0020            
						   33727 => x"20",
						   33728 => x"44",		-- 0083c0: 449C            
						   33729 => x"9C",
						   33730 => x"34",		-- 0083c2: 3440             MOV.W   #0x2000,R4
						   33731 => x"60",
						   33732 => x"00",		-- 0083c4: 0020            
						   33733 => x"20",
						   33734 => x"90",		-- 0083c6: 9010             SWPB    Var1
						   33735 => x"30",
						   33736 => x"3C",		-- 0083c8: 3C9C            
						   33737 => x"9C",
						   33738 => x"94",		-- 0083ca: 9410             SWPB    0x0004(R4)
						   33739 => x"30",
						   33740 => x"04",		-- 0083cc: 0400            
						   33741 => x"00",
						   33742 => x"34",		-- 0083ce: 3440             MOV.W   #0x00ff,R4
						   33743 => x"60",
						   33744 => x"FF",		-- 0083d0: FF00            
						   33745 => x"00",
						   33746 => x"84",		-- 0083d2: 8411             SXT     R4
						   33747 => x"31",
						   33748 => x"90",		-- 0083d4: 9011             SXT     Const2
						   33749 => x"31",
						   33750 => x"4C",		-- 0083d6: 4C9C            
						   33751 => x"9C",
						   33752 => x"92",		-- 0083d8: 9211             SXT     &Con1
						   33753 => x"31",
						   33754 => x"00",		-- 0083da: 0020            
						   33755 => x"20",
						   33756 => x"B0",		-- 0083dc: B040             MOV.W   #0x2000,Var1
						   33757 => x"60",
						   33758 => x"00",		-- 0083de: 0020            
						   33759 => x"20",
						   33760 => x"24",		-- 0083e0: 249C            
						   33761 => x"9C",
						   33762 => x"34",		-- 0083e2: 3440             MOV.W   #0x2000,R4
						   33763 => x"60",
						   33764 => x"00",		-- 0083e4: 0020            
						   33765 => x"20",
						   33766 => x"90",		-- 0083e6: 9011             SXT     Var1
						   33767 => x"31",
						   33768 => x"1C",		-- 0083e8: 1C9C            
						   33769 => x"9C",
						   33770 => x"94",		-- 0083ea: 9411             SXT     0x0004(R4)
						   33771 => x"31",
						   33772 => x"04",		-- 0083ec: 0400            
						   33773 => x"00",
						   33774 => x"12",		-- 0083ee: 12D3             SETC    
						   33775 => x"F3",
						   33776 => x"22",		-- 0083f0: 22D2             SETN    
						   33777 => x"F2",
						   33778 => x"22",		-- 0083f2: 22D3             SETZ    
						   33779 => x"F3",
						   33780 => x"12",		-- 0083f4: 12C3             CLRC    
						   33781 => x"E3",
						   33782 => x"22",		-- 0083f6: 22C2             CLRN    
						   33783 => x"E2",
						   33784 => x"22",		-- 0083f8: 22C3             CLRZ    
						   33785 => x"E3",
						   33786 => x"3A",		-- 0083fa: 3A40             MOV.W   #0x001c,R10
						   33787 => x"60",
						   33788 => x"1C",		-- 0083fc: 1C00            
						   33789 => x"00",
						   33790 => x"0A",		-- 0083fe: 0A43             CLR.W   R10
						   33791 => x"63",
						   33792 => x"80",		-- 008400: 8043             CLR.W   Var1
						   33793 => x"63",
						   33794 => x"02",		-- 008402: 029C            
						   33795 => x"9C",
						   33796 => x"82",		-- 008404: 8243             CLR.W   &Con1
						   33797 => x"63",
						   33798 => x"00",		-- 008406: 0020            
						   33799 => x"20",
						   33800 => x"3A",		-- 008408: 3A40             MOV.W   #0x2000,R10
						   33801 => x"60",
						   33802 => x"00",		-- 00840a: 0020            
						   33803 => x"20",
						   33804 => x"8A",		-- 00840c: 8A43             CLR.W   0x0002(R10)
						   33805 => x"63",
						   33806 => x"02",		-- 00840e: 0200            
						   33807 => x"00",
						   33808 => x"12",		-- 008410: 12D3             SETC    
						   33809 => x"F3",
						   33810 => x"00",		-- 008412: 002C             JHS     (_jc)
						   33811 => x"4C",
						   33812 => x"12",		-- 008414: 12C3             CLRC    
						   33813 => x"E3",
						   33814 => x"FE",		-- 008416: FE2F             JHS     (_jc)
						   33815 => x"4F",
						   33816 => x"12",		-- 008418: 12D3             SETC    
						   33817 => x"F3",
						   33818 => x"00",		-- 00841a: 002C             JHS     (_jhs)
						   33819 => x"4C",
						   33820 => x"12",		-- 00841c: 12C3             CLRC    
						   33821 => x"E3",
						   33822 => x"FE",		-- 00841e: FE2F             JHS     (_jhs)
						   33823 => x"4F",
						   33824 => x"22",		-- 008420: 22D3             SETZ    
						   33825 => x"F3",
						   33826 => x"00",		-- 008422: 0024             JEQ     (_jeq)
						   33827 => x"44",
						   33828 => x"22",		-- 008424: 22C3             CLRZ    
						   33829 => x"E3",
						   33830 => x"FE",		-- 008426: FE27             JEQ     (_jeq)
						   33831 => x"47",
						   33832 => x"22",		-- 008428: 22D3             SETZ    
						   33833 => x"F3",
						   33834 => x"00",		-- 00842a: 0024             JEQ     (_jz)
						   33835 => x"44",
						   33836 => x"22",		-- 00842c: 22C3             CLRZ    
						   33837 => x"E3",
						   33838 => x"FE",		-- 00842e: FE27             JEQ     (_jz)
						   33839 => x"47",
						   33840 => x"14",		-- 008430: 1443             MOV.W   #1,R4
						   33841 => x"63",
						   33842 => x"04",		-- 008432: 0493             TST.W   R4
						   33843 => x"B3",
						   33844 => x"00",		-- 008434: 0034             JGE     (_jge)
						   33845 => x"54",
						   33846 => x"04",		-- 008436: 0443             CLR.W   R4
						   33847 => x"63",
						   33848 => x"14",		-- 008438: 1493             CMP.W   #1,R4
						   33849 => x"B3",
						   33850 => x"FD",		-- 00843a: FD37             JGE     (_jge)
						   33851 => x"57",
						   33852 => x"04",		-- 00843c: 0443             CLR.W   R4
						   33853 => x"63",
						   33854 => x"14",		-- 00843e: 1493             CMP.W   #1,R4
						   33855 => x"B3",
						   33856 => x"00",		-- 008440: 0038             JL      (_jl)
						   33857 => x"58",
						   33858 => x"14",		-- 008442: 1443             MOV.W   #1,R4
						   33859 => x"63",
						   33860 => x"04",		-- 008444: 0493             TST.W   R4
						   33861 => x"B3",
						   33862 => x"FD",		-- 008446: FD3B             JL      (_jl)
						   33863 => x"5B",
						   33864 => x"00",		-- 008448: 003C             JMP     (_jmp)
						   33865 => x"5C",
						   33866 => x"03",		-- 00844a: 0343             NOP     
						   33867 => x"63",
						   33868 => x"22",		-- 00844c: 22D2             SETN    
						   33869 => x"F2",
						   33870 => x"00",		-- 00844e: 0030             JN      (_jn)
						   33871 => x"50",
						   33872 => x"22",		-- 008450: 22C2             CLRN    
						   33873 => x"E2",
						   33874 => x"FE",		-- 008452: FE33             JN      (_jn)
						   33875 => x"53",
						   33876 => x"22",		-- 008454: 22C2             CLRN    
						   33877 => x"E2",
						   33878 => x"00",		-- 008456: 0028             JLO     (_jnc)
						   33879 => x"48",
						   33880 => x"22",		-- 008458: 22D2             SETN    
						   33881 => x"F2",
						   33882 => x"FE",		-- 00845a: FE2B             JLO     (_jnc)
						   33883 => x"4B",
						   33884 => x"22",		-- 00845c: 22C2             CLRN    
						   33885 => x"E2",
						   33886 => x"00",		-- 00845e: 0028             JLO     (_jlo)
						   33887 => x"48",
						   33888 => x"22",		-- 008460: 22D2             SETN    
						   33889 => x"F2",
						   33890 => x"FE",		-- 008462: FE2B             JLO     (_jlo)
						   33891 => x"4B",
						   33892 => x"22",		-- 008464: 22C3             CLRZ    
						   33893 => x"E3",
						   33894 => x"00",		-- 008466: 0020             JNE     (_jne)
						   33895 => x"40",
						   33896 => x"22",		-- 008468: 22D3             SETZ    
						   33897 => x"F3",
						   33898 => x"FE",		-- 00846a: FE23             JNE     (_jne)
						   33899 => x"43",
						   33900 => x"22",		-- 00846c: 22C3             CLRZ    
						   33901 => x"E3",
						   33902 => x"00",		-- 00846e: 0020             JNE     (_jnz)
						   33903 => x"40",
						   33904 => x"22",		-- 008470: 22D3             SETZ    
						   33905 => x"F3",
						   33906 => x"FE",		-- 008472: FE23             JNE     (_jnz)
						   33907 => x"43",
						   33908 => x"34",		-- 008474: 3440             MOV.W   #0x847a,R4
						   33909 => x"60",
						   33910 => x"7A",		-- 008476: 7A84            
						   33911 => x"84",
						   33912 => x"00",		-- 008478: 0044             BR      R4
						   33913 => x"64",
						   33914 => x"B0",		-- 00847a: B040             MOV.W   #0x8484,Const2
						   33915 => x"60",
						   33916 => x"84",		-- 00847c: 8484            
						   33917 => x"84",
						   33918 => x"A4",		-- 00847e: A49B            
						   33919 => x"9B",
						   33920 => x"10",		-- 008480: 1040             BR      Const2
						   33921 => x"60",
						   33922 => x"A0",		-- 008482: A09B            
						   33923 => x"9B",
						   33924 => x"30",		-- 008484: 3040             BR      #br_3
						   33925 => x"60",
						   33926 => x"88",		-- 008486: 8884            
						   33927 => x"84",
						   33928 => x"03",		-- 008488: 0343             NOP     
						   33929 => x"63",
						   33930 => x"34",		-- 00848a: 3440             MOV.W   #0x00ff,R4
						   33931 => x"60",
						   33932 => x"FF",		-- 00848c: FF00            
						   33933 => x"00",
						   33934 => x"30",		-- 00848e: 3012             PUSH    #0xf0f0
						   33935 => x"32",
						   33936 => x"F0",		-- 008490: F0F0            
						   33937 => x"F0",
						   33938 => x"04",		-- 008492: 0412             PUSH    R4
						   33939 => x"32",
						   33940 => x"12",		-- 008494: 1212             PUSH    &Con1
						   33941 => x"32",
						   33942 => x"00",		-- 008496: 0020            
						   33943 => x"20",
						   33944 => x"34",		-- 008498: 3440             MOV.W   #0x2000,R4
						   33945 => x"60",
						   33946 => x"00",		-- 00849a: 0020            
						   33947 => x"20",
						   33948 => x"14",		-- 00849c: 1412             PUSH    0x0000(R4)
						   33949 => x"32",
						   33950 => x"00",		-- 00849e: 0000            
						   33951 => x"00",
						   33952 => x"30",		-- 0084a0: 3012             PUSH    #0x2000
						   33953 => x"32",
						   33954 => x"00",		-- 0084a2: 0020            
						   33955 => x"20",
						   33956 => x"35",		-- 0084a4: 3512             PUSH    @R5+
						   33957 => x"32",
						   33958 => x"34",		-- 0084a6: 3441             POP.W   R4
						   33959 => x"61",
						   33960 => x"B0",		-- 0084a8: B041             POP.W   Const2
						   33961 => x"61",
						   33962 => x"78",		-- 0084aa: 789B            
						   33963 => x"9B",
						   33964 => x"B2",		-- 0084ac: B241             POP.W   &Con1
						   33965 => x"61",
						   33966 => x"00",		-- 0084ae: 0020            
						   33967 => x"20",
						   33968 => x"B0",		-- 0084b0: B040             MOV.W   #0x2000,Var1
						   33969 => x"60",
						   33970 => x"00",		-- 0084b2: 0020            
						   33971 => x"20",
						   33972 => x"50",		-- 0084b4: 509B            
						   33973 => x"9B",
						   33974 => x"34",		-- 0084b6: 3440             MOV.W   #0x2000,R4
						   33975 => x"60",
						   33976 => x"00",		-- 0084b8: 0020            
						   33977 => x"20",
						   33978 => x"B0",		-- 0084ba: B041             POP.W   Var1
						   33979 => x"61",
						   33980 => x"48",		-- 0084bc: 489B            
						   33981 => x"9B",
						   33982 => x"B4",		-- 0084be: B441             POP.W   0x0004(R4)
						   33983 => x"61",
						   33984 => x"04",		-- 0084c0: 0400            
						   33985 => x"00",
						   33986 => x"34",		-- 0084c2: 3441             POP.W   R4
						   33987 => x"61",
						   33988 => x"05",		-- 0084c4: 0543             CLR.W   R5
						   33989 => x"63",
						   33990 => x"34",		-- 0084c6: 3440             MOV.W   #0x84e4,R4
						   33991 => x"60",
						   33992 => x"E4",		-- 0084c8: E484            
						   33993 => x"84",
						   33994 => x"B0",		-- 0084ca: B040             MOV.W   #0x84e4,Var1
						   33995 => x"60",
						   33996 => x"E4",		-- 0084cc: E484            
						   33997 => x"84",
						   33998 => x"36",		-- 0084ce: 369B            
						   33999 => x"9B",
						   34000 => x"B0",		-- 0084d0: B012             CALL    #add_3
						   34001 => x"32",
						   34002 => x"E4",		-- 0084d2: E484            
						   34003 => x"84",
						   34004 => x"84",		-- 0084d4: 8412             CALL    R4
						   34005 => x"32",
						   34006 => x"90",		-- 0084d6: 9012             CALL    Var1
						   34007 => x"32",
						   34008 => x"2C",		-- 0084d8: 2C9B            
						   34009 => x"9B",
						   34010 => x"B0",		-- 0084da: B012             CALL    #add_3
						   34011 => x"32",
						   34012 => x"E4",		-- 0084dc: E484            
						   34013 => x"84",
						   34014 => x"30",		-- 0084de: 3040             BR      #main
						   34015 => x"60",
						   34016 => x"3E",		-- 0084e0: 3E80            
						   34017 => x"80",
						   34018 => x"03",		-- 0084e2: 0343             NOP     
						   34019 => x"63",
						   34020 => x"35",		-- 0084e4: 3550             ADD.W   #0x0003,R5
						   34021 => x"70",
						   34022 => x"03",		-- 0084e6: 0300            
						   34023 => x"00",
						   34024 => x"30",		-- 0084e8: 3041             RET     
						   34025 => x"61",
						   34026 => x"32",		-- 0084ea: 32D0             BIS.W   #0x0010,SR
						   34027 => x"F0",
        -- IRQ Vectors (Interrupts)
                           65534 =>  x"00",		-- Reset Vector = xFFFE:xFFFF
                           65535 =>  x"80",		--  Startup Value = x8000

                           others => x"00");

    signal EN : std_logic;

    begin
    -- Note 1:  The bus system uses a 16-bit Address (MAB)
    --          This address size can access locations from x0000 to xFFFF
    --          But our array is only defined from x8000 to xFFFF and
    --          if we try to access it with any other address, it will crash.
    --          So the first thing we need to do is create a local enable that
    --          will only assert when MAB is within x8000 to xFFFF.

     LOCAL_EN : process (MAB) 
       begin
         if ( (to_integer(unsigned(MAB)) >= 32768) and (to_integer(unsigned(MAB)) <= 65535)) then
           EN <= '1';
         else 
           EN <= '0';
        end if;
      end process;


    -- Note 2:  The bus system uses a 16-bit Address (MAB)
    --          The MDB_out is also provided as a 16-bit word
    --          However, the memory array is actually built as 8-bit bytes.
    --          So for a given 16-bit MAB, we give MDB_out = HB : LB
    --                                                 or  = ROM(MAB);1) : ROM(MAB)

    MEMORY_ROM : process (clk) 
     begin
        if (rising_edge(clk)) then
            if (EN='1' and write='0') then                      
              MDB_in <= ROM(to_integer(unsigned(MAB)) + 1 ) & ROM(to_integer(unsigned(MAB))); 
            end if;
      end if;
   end process;


end architecture;