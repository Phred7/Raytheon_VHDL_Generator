library IEEE;
    use IEEE.std_logic_1164.all;
    use IEEE.numeric_std.all;
    package highroller is
    constant FORMAT_2 : integer := 3;
    constant JMP1 : integer := 4;
    constant JMP2 : integer := 5;
    constant MOV : integer := 6;
    constant OFFSET : integer := 2;
    end highroller;
