library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;


entity highroller_memory is
    port ( clk	: in	std_logic;
         MAB		: in	std_logic_vector(15 downto 0);
         MDB_in  	: out	std_logic_vector(15 downto 0);
         MDB_out  	: in	std_logic_vector(15 downto 0);
         write	    : in	std_logic);
end entity;

architecture highroller_memory_arch of highroller_memory is

type rom_type is array (32768 to 65535) of std_logic_vector(7 downto 0);  -- this is MAB: x8000 to xFFFF
    
constant ROM : rom_type :=(32768 => x"31",		-- 008000: 3140             MOV.W   #0x3000,SP
						   32769 => x"60",
						   32770 => x"00",		-- 008002: 0030            
						   32771 => x"30",
						   32772 => x"B2",		-- 008004: B240             MOV.W   #0x5a80,&WDTCTL_L
						   32773 => x"60",
						   32774 => x"80",		-- 008006: 805A            
						   32775 => x"5A",
						   32776 => x"CC",		-- 008008: CC01            
						   32777 => x"01",
						   32778 => x"34",		-- 00800a: 3440             MOV.W   #0x2000,R4
						   32779 => x"60",
						   32780 => x"00",		-- 00800c: 0020            
						   32781 => x"20",
						   32782 => x"05",		-- 00800e: 0544             MOV.W   R4,R5
						   32783 => x"64",
						   32784 => x"36",		-- 008010: 3640             MOV.W   #0x2004,R6
						   32785 => x"60",
						   32786 => x"04",		-- 008012: 0420            
						   32787 => x"20",
						   32788 => x"E2",		-- 008014: E2C3             BIC.B   #2,&P4DIR
						   32789 => x"E3",
						   32790 => x"25",		-- 008016: 2502            
						   32791 => x"02",
						   32792 => x"E2",		-- 008018: E2D3             BIS.B   #2,&P4REN
						   32793 => x"F3",
						   32794 => x"27",		-- 00801a: 2702            
						   32795 => x"02",
						   32796 => x"E2",		-- 00801c: E2D3             BIS.B   #2,&P4OUT
						   32797 => x"F3",
						   32798 => x"23",		-- 00801e: 2302            
						   32799 => x"02",
						   32800 => x"F2",		-- 008020: F2C3             BIC.B   #-1,&P4IFG
						   32801 => x"E3",
						   32802 => x"3D",		-- 008022: 3D02            
						   32803 => x"02",
						   32804 => x"E2",		-- 008024: E2D3             BIS.B   #2,&P4IES
						   32805 => x"F3",
						   32806 => x"39",		-- 008026: 3902            
						   32807 => x"02",
						   32808 => x"E2",		-- 008028: E2D3             BIS.B   #2,&P4IE
						   32809 => x"F3",
						   32810 => x"3B",		-- 00802a: 3B02            
						   32811 => x"02",
						   32812 => x"03",		-- 00802c: 0343             NOP     
						   32813 => x"63",
						   32814 => x"03",		-- 008030: 0343             NOP     
						   32815 => x"63",
						   32816 => x"03",		-- 008034: 0343             NOP     
						   32817 => x"63",
						   32818 => x"03",		-- 008038: 0343             NOP     
						   32819 => x"63",
						   32820 => x"D2",		-- 00803a: D2C3             BIC.B   #1,&PM5CTL0_L
						   32821 => x"E3",
						   32822 => x"30",		-- 00803c: 3001            
						   32823 => x"01",
						   32824 => x"17",		-- 00803e: 1742             MOV.W   &Con1,R7
						   32825 => x"62",
						   32826 => x"00",		-- 008040: 0020            
						   32827 => x"20",
						   32828 => x"18",		-- 008042: 1840             MOV.W   Con2,R8
						   32829 => x"60",
						   32830 => x"BE",		-- 008044: BE9F            
						   32831 => x"9F",
						   32832 => x"29",		-- 008046: 2944             MOV.W   @R4,R9
						   32833 => x"64",
						   32834 => x"3A",		-- 008048: 3A45             MOV.W   @R5+,R10
						   32835 => x"65",
						   32836 => x"3B",		-- 00804a: 3B45             MOV.W   @R5+,R11
						   32837 => x"65",
						   32838 => x"96",		-- 00804c: 9644             MOV.W   0x0002(R4),0x0004(R6)
						   32839 => x"64",
						   32840 => x"02",		-- 00804e: 0200            
						   32841 => x"00",
						   32842 => x"04",		-- 008050: 0400            
						   32843 => x"00",
						   32844 => x"34",		-- 008052: 3440             MOV.W   #0x2000,R4
						   32845 => x"60",
						   32846 => x"00",		-- 008054: 0020            
						   32847 => x"20",
						   32848 => x"80",		-- 008056: 8054             ADD.W   R4,Const2
						   32849 => x"74",
						   32850 => x"CA",		-- 008058: CA9F            
						   32851 => x"9F",
						   32852 => x"15",		-- 00805a: 1552             ADD.W   &Con1,R5
						   32853 => x"72",
						   32854 => x"00",		-- 00805c: 0020            
						   32855 => x"20",
						   32856 => x"34",		-- 00805e: 3440             MOV.W   #0x2000,R4
						   32857 => x"60",
						   32858 => x"00",		-- 008060: 0020            
						   32859 => x"20",
						   32860 => x"36",		-- 008062: 3640             MOV.W   #0x2004,R6
						   32861 => x"60",
						   32862 => x"04",		-- 008064: 0420            
						   32863 => x"20",
						   32864 => x"A6",		-- 008066: A654             ADD.W   @R4,0x0004(R6)
						   32865 => x"74",
						   32866 => x"04",		-- 008068: 0400            
						   32867 => x"00",
						   32868 => x"B0",		-- 00806a: B050             ADD.W   #0x2000,Var1
						   32869 => x"70",
						   32870 => x"00",		-- 00806c: 0020            
						   32871 => x"20",
						   32872 => x"96",		-- 00806e: 969F            
						   32873 => x"9F",
						   32874 => x"36",		-- 008070: 3655             ADD.W   @R5+,R6
						   32875 => x"75",
						   32876 => x"05",		-- 008072: 0564             ADDC.W  R4,R5
						   32877 => x"84",
						   32878 => x"80",		-- 008074: 8065             ADDC.W  R5,Const2
						   32879 => x"85",
						   32880 => x"AC",		-- 008076: AC9F            
						   32881 => x"9F",
						   32882 => x"15",		-- 008078: 1562             ADDC.W  &Con1,R5
						   32883 => x"82",
						   32884 => x"00",		-- 00807a: 0020            
						   32885 => x"20",
						   32886 => x"34",		-- 00807c: 3440             MOV.W   #0x2000,R4
						   32887 => x"60",
						   32888 => x"00",		-- 00807e: 0020            
						   32889 => x"20",
						   32890 => x"36",		-- 008080: 3640             MOV.W   #0x2004,R6
						   32891 => x"60",
						   32892 => x"04",		-- 008082: 0420            
						   32893 => x"20",
						   32894 => x"A6",		-- 008084: A664             ADDC.W  @R4,0x0004(R6)
						   32895 => x"84",
						   32896 => x"04",		-- 008086: 0400            
						   32897 => x"00",
						   32898 => x"B0",		-- 008088: B060             ADDC.W  #0x2000,Var1
						   32899 => x"80",
						   32900 => x"00",		-- 00808a: 0020            
						   32901 => x"20",
						   32902 => x"78",		-- 00808c: 789F            
						   32903 => x"9F",
						   32904 => x"36",		-- 00808e: 3665             ADDC.W  @R5+,R6
						   32905 => x"85",
						   32906 => x"04",		-- 008092: 0463             ADC.W   R4
						   32907 => x"83",
						   32908 => x"80",		-- 008094: 8063             ADC.W   Const2
						   32909 => x"83",
						   32910 => x"8C",		-- 008096: 8C9F            
						   32911 => x"9F",
						   32912 => x"82",		-- 008098: 8263             ADC.W   &Con1
						   32913 => x"83",
						   32914 => x"00",		-- 00809a: 0020            
						   32915 => x"20",
						   32916 => x"B0",		-- 00809c: B040             MOV.W   #0x2000,Var1
						   32917 => x"60",
						   32918 => x"00",		-- 00809e: 0020            
						   32919 => x"20",
						   32920 => x"64",		-- 0080a0: 649F            
						   32921 => x"9F",
						   32922 => x"34",		-- 0080a2: 3440             MOV.W   #0x2000,R4
						   32923 => x"60",
						   32924 => x"00",		-- 0080a4: 0020            
						   32925 => x"20",
						   32926 => x"80",		-- 0080a8: 8063             ADC.W   Var1
						   32927 => x"83",
						   32928 => x"5A",		-- 0080aa: 5A9F            
						   32929 => x"9F",
						   32930 => x"84",		-- 0080ac: 8463             ADC.W   0x0004(R4)
						   32931 => x"83",
						   32932 => x"04",		-- 0080ae: 0400            
						   32933 => x"00",
						   32934 => x"05",		-- 0080b0: 0584             SUB.W   R4,R5
						   32935 => x"A4",
						   32936 => x"80",		-- 0080b2: 8084             SUB.W   R4,Const2
						   32937 => x"A4",
						   32938 => x"6E",		-- 0080b4: 6E9F            
						   32939 => x"9F",
						   32940 => x"15",		-- 0080b6: 1582             SUB.W   &Con1,R5
						   32941 => x"A2",
						   32942 => x"00",		-- 0080b8: 0020            
						   32943 => x"20",
						   32944 => x"34",		-- 0080ba: 3440             MOV.W   #0x2000,R4
						   32945 => x"60",
						   32946 => x"00",		-- 0080bc: 0020            
						   32947 => x"20",
						   32948 => x"36",		-- 0080be: 3640             MOV.W   #0x2004,R6
						   32949 => x"60",
						   32950 => x"04",		-- 0080c0: 0420            
						   32951 => x"20",
						   32952 => x"A6",		-- 0080c2: A684             SUB.W   @R4,0x0004(R6)
						   32953 => x"A4",
						   32954 => x"04",		-- 0080c4: 0400            
						   32955 => x"00",
						   32956 => x"B0",		-- 0080c6: B080             SUB.W   #0x2000,Var1
						   32957 => x"A0",
						   32958 => x"00",		-- 0080c8: 0020            
						   32959 => x"20",
						   32960 => x"3A",		-- 0080ca: 3A9F            
						   32961 => x"9F",
						   32962 => x"36",		-- 0080cc: 3685             SUB.W   @R5+,R6
						   32963 => x"A5",
						   32964 => x"06",		-- 0080ce: 0675             SUBC.W  R5,R6
						   32965 => x"95",
						   32966 => x"80",		-- 0080d0: 8074             SUBC.W  R4,Const2
						   32967 => x"94",
						   32968 => x"50",		-- 0080d2: 509F            
						   32969 => x"9F",
						   32970 => x"15",		-- 0080d4: 1572             SUBC.W  &Con1,R5
						   32971 => x"92",
						   32972 => x"00",		-- 0080d6: 0020            
						   32973 => x"20",
						   32974 => x"34",		-- 0080d8: 3440             MOV.W   #0x2000,R4
						   32975 => x"60",
						   32976 => x"00",		-- 0080da: 0020            
						   32977 => x"20",
						   32978 => x"36",		-- 0080dc: 3640             MOV.W   #0x2004,R6
						   32979 => x"60",
						   32980 => x"04",		-- 0080de: 0420            
						   32981 => x"20",
						   32982 => x"A6",		-- 0080e0: A674             SUBC.W  @R4,0x0004(R6)
						   32983 => x"94",
						   32984 => x"04",		-- 0080e2: 0400            
						   32985 => x"00",
						   32986 => x"B0",		-- 0080e4: B070             SUBC.W  #0x2000,Var1
						   32987 => x"90",
						   32988 => x"00",		-- 0080e6: 0020            
						   32989 => x"20",
						   32990 => x"1C",		-- 0080e8: 1C9F            
						   32991 => x"9F",
						   32992 => x"36",		-- 0080ea: 3675             SUBC.W  @R5+,R6
						   32993 => x"95",
						   32994 => x"30",		-- 0080f2: 309F            
						   32995 => x"9F",
						   32996 => x"00",		-- 0080f6: 0020            
						   32997 => x"20",
						   32998 => x"B0",		-- 0080f8: B040             MOV.W   #0x2000,Var1
						   32999 => x"60",
						   33000 => x"00",		-- 0080fa: 0020            
						   33001 => x"20",
						   33002 => x"08",		-- 0080fc: 089F            
						   33003 => x"9F",
						   33004 => x"34",		-- 0080fe: 3440             MOV.W   #0x2000,R4
						   33005 => x"60",
						   33006 => x"00",		-- 008100: 0020            
						   33007 => x"20",
						   33008 => x"FE",		-- 008106: FE9E            
						   33009 => x"9E",
						   33010 => x"04",		-- 00810a: 0400            
						   33011 => x"00",
						   33012 => x"05",		-- 00810e: 05A4             DADD.W  R4,R5
						   33013 => x"C4",
						   33014 => x"80",		-- 008110: 80A4             DADD.W  R4,Const2
						   33015 => x"C4",
						   33016 => x"10",		-- 008112: 109F            
						   33017 => x"9F",
						   33018 => x"15",		-- 008114: 15A2             DADD.W  &Con1,R5
						   33019 => x"C2",
						   33020 => x"00",		-- 008116: 0020            
						   33021 => x"20",
						   33022 => x"34",		-- 008118: 3440             MOV.W   #0x2000,R4
						   33023 => x"60",
						   33024 => x"00",		-- 00811a: 0020            
						   33025 => x"20",
						   33026 => x"36",		-- 00811c: 3640             MOV.W   #0x2004,R6
						   33027 => x"60",
						   33028 => x"04",		-- 00811e: 0420            
						   33029 => x"20",
						   33030 => x"A6",		-- 008122: A6A4             DADD.W  @R4,0x0004(R6)
						   33031 => x"C4",
						   33032 => x"04",		-- 008124: 0400            
						   33033 => x"00",
						   33034 => x"B0",		-- 008126: B0A0             DADD.W  #0x2000,Var1
						   33035 => x"C0",
						   33036 => x"00",		-- 008128: 0020            
						   33037 => x"20",
						   33038 => x"DA",		-- 00812a: DA9E            
						   33039 => x"9E",
						   33040 => x"36",		-- 00812c: 36A5             DADD.W  @R5+,R6
						   33041 => x"C5",
						   33042 => x"04",		-- 008130: 04A3             DADC.W  R4
						   33043 => x"C3",
						   33044 => x"80",		-- 008132: 80A3             DADC.W  Const2
						   33045 => x"C3",
						   33046 => x"EE",		-- 008134: EE9E            
						   33047 => x"9E",
						   33048 => x"82",		-- 008136: 82A3             DADC.W  &Con1
						   33049 => x"C3",
						   33050 => x"00",		-- 008138: 0020            
						   33051 => x"20",
						   33052 => x"B0",		-- 00813a: B040             MOV.W   #0x2000,Var1
						   33053 => x"60",
						   33054 => x"00",		-- 00813c: 0020            
						   33055 => x"20",
						   33056 => x"C6",		-- 00813e: C69E            
						   33057 => x"9E",
						   33058 => x"34",		-- 008140: 3440             MOV.W   #0x2000,R4
						   33059 => x"60",
						   33060 => x"00",		-- 008142: 0020            
						   33061 => x"20",
						   33062 => x"80",		-- 008146: 80A3             DADC.W  Var1
						   33063 => x"C3",
						   33064 => x"BC",		-- 008148: BC9E            
						   33065 => x"9E",
						   33066 => x"84",		-- 00814a: 84A3             DADC.W  0x0004(R4)
						   33067 => x"C3",
						   33068 => x"04",		-- 00814c: 0400            
						   33069 => x"00",
						   33070 => x"14",		-- 00814e: 1453             INC.W   R4
						   33071 => x"73",
						   33072 => x"90",		-- 008150: 9053             INC.W   Const2
						   33073 => x"73",
						   33074 => x"D0",		-- 008152: D09E            
						   33075 => x"9E",
						   33076 => x"92",		-- 008154: 9253             INC.W   &Con1
						   33077 => x"73",
						   33078 => x"00",		-- 008156: 0020            
						   33079 => x"20",
						   33080 => x"B0",		-- 008158: B040             MOV.W   #0x2000,Var1
						   33081 => x"60",
						   33082 => x"00",		-- 00815a: 0020            
						   33083 => x"20",
						   33084 => x"A8",		-- 00815c: A89E            
						   33085 => x"9E",
						   33086 => x"34",		-- 00815e: 3440             MOV.W   #0x2000,R4
						   33087 => x"60",
						   33088 => x"00",		-- 008160: 0020            
						   33089 => x"20",
						   33090 => x"90",		-- 008162: 9053             INC.W   Var1
						   33091 => x"73",
						   33092 => x"A0",		-- 008164: A09E            
						   33093 => x"9E",
						   33094 => x"94",		-- 008166: 9453             INC.W   0x0004(R4)
						   33095 => x"73",
						   33096 => x"04",		-- 008168: 0400            
						   33097 => x"00",
						   33098 => x"24",		-- 00816a: 2453             INCD.W  R4
						   33099 => x"73",
						   33100 => x"A0",		-- 00816c: A053             INCD.W  Const2
						   33101 => x"73",
						   33102 => x"B4",		-- 00816e: B49E            
						   33103 => x"9E",
						   33104 => x"A2",		-- 008170: A253             INCD.W  &Con1
						   33105 => x"73",
						   33106 => x"00",		-- 008172: 0020            
						   33107 => x"20",
						   33108 => x"B0",		-- 008174: B040             MOV.W   #0x2000,Var1
						   33109 => x"60",
						   33110 => x"00",		-- 008176: 0020            
						   33111 => x"20",
						   33112 => x"8C",		-- 008178: 8C9E            
						   33113 => x"9E",
						   33114 => x"34",		-- 00817a: 3440             MOV.W   #0x2000,R4
						   33115 => x"60",
						   33116 => x"00",		-- 00817c: 0020            
						   33117 => x"20",
						   33118 => x"A0",		-- 00817e: A053             INCD.W  Var1
						   33119 => x"73",
						   33120 => x"84",		-- 008180: 849E            
						   33121 => x"9E",
						   33122 => x"A4",		-- 008182: A453             INCD.W  0x0004(R4)
						   33123 => x"73",
						   33124 => x"04",		-- 008184: 0400            
						   33125 => x"00",
						   33126 => x"14",		-- 008186: 1483             DEC.W   R4
						   33127 => x"A3",
						   33128 => x"90",		-- 008188: 9083             DEC.W   Const2
						   33129 => x"A3",
						   33130 => x"98",		-- 00818a: 989E            
						   33131 => x"9E",
						   33132 => x"92",		-- 00818c: 9283             DEC.W   &Con1
						   33133 => x"A3",
						   33134 => x"00",		-- 00818e: 0020            
						   33135 => x"20",
						   33136 => x"B0",		-- 008190: B040             MOV.W   #0x2000,Var1
						   33137 => x"60",
						   33138 => x"00",		-- 008192: 0020            
						   33139 => x"20",
						   33140 => x"70",		-- 008194: 709E            
						   33141 => x"9E",
						   33142 => x"34",		-- 008196: 3440             MOV.W   #0x2000,R4
						   33143 => x"60",
						   33144 => x"00",		-- 008198: 0020            
						   33145 => x"20",
						   33146 => x"90",		-- 00819a: 9083             DEC.W   Var1
						   33147 => x"A3",
						   33148 => x"68",		-- 00819c: 689E            
						   33149 => x"9E",
						   33150 => x"94",		-- 00819e: 9483             DEC.W   0x0004(R4)
						   33151 => x"A3",
						   33152 => x"04",		-- 0081a0: 0400            
						   33153 => x"00",
						   33154 => x"24",		-- 0081a2: 2483             DECD.W  R4
						   33155 => x"A3",
						   33156 => x"A0",		-- 0081a4: A083             DECD.W  Const2
						   33157 => x"A3",
						   33158 => x"7C",		-- 0081a6: 7C9E            
						   33159 => x"9E",
						   33160 => x"A2",		-- 0081a8: A283             DECD.W  &Con1
						   33161 => x"A3",
						   33162 => x"00",		-- 0081aa: 0020            
						   33163 => x"20",
						   33164 => x"B0",		-- 0081ac: B040             MOV.W   #0x2000,Var1
						   33165 => x"60",
						   33166 => x"00",		-- 0081ae: 0020            
						   33167 => x"20",
						   33168 => x"54",		-- 0081b0: 549E            
						   33169 => x"9E",
						   33170 => x"34",		-- 0081b2: 3440             MOV.W   #0x2000,R4
						   33171 => x"60",
						   33172 => x"00",		-- 0081b4: 0020            
						   33173 => x"20",
						   33174 => x"A0",		-- 0081b6: A083             DECD.W  Var1
						   33175 => x"A3",
						   33176 => x"4C",		-- 0081b8: 4C9E            
						   33177 => x"9E",
						   33178 => x"A4",		-- 0081ba: A483             DECD.W  0x0004(R4)
						   33179 => x"A3",
						   33180 => x"04",		-- 0081bc: 0400            
						   33181 => x"00",
						   33182 => x"74",		-- 0081be: 7440             MOV.B   #0x004e,R4
						   33183 => x"60",
						   33184 => x"4E",		-- 0081c0: 4E00            
						   33185 => x"00",
						   33186 => x"34",		-- 0081c4: 3440             MOV.W   #0x2032,R4
						   33187 => x"60",
						   33188 => x"32",		-- 0081c6: 3220            
						   33189 => x"20",
						   33190 => x"20",		-- 0081cc: 2020            
						   33191 => x"20",
						   33192 => x"62",		-- 0081d0: 629E            
						   33193 => x"9E",
						   33194 => x"34",		-- 0081d2: 3440             MOV.W   #0x2032,R4
						   33195 => x"60",
						   33196 => x"32",		-- 0081d4: 3220            
						   33197 => x"20",
						   33198 => x"02",		-- 0081d8: 0200            
						   33199 => x"00",
						   33200 => x"74",		-- 0081da: 7440             MOV.B   #0x00aa,R4
						   33201 => x"60",
						   33202 => x"AA",		-- 0081dc: AA00            
						   33203 => x"00",
						   33204 => x"74",		-- 0081de: 74F0             AND.B   #0x000f,R4
						   33205 => x"10",
						   33206 => x"0F",		-- 0081e0: 0F00            
						   33207 => x"00",
						   33208 => x"05",		-- 0081e2: 05F4             AND.W   R4,R5
						   33209 => x"14",
						   33210 => x"80",		-- 0081e4: 80F4             AND.W   R4,Const2
						   33211 => x"14",
						   33212 => x"3C",		-- 0081e6: 3C9E            
						   33213 => x"9E",
						   33214 => x"15",		-- 0081e8: 15F2             AND.W   &Con1,R5
						   33215 => x"12",
						   33216 => x"00",		-- 0081ea: 0020            
						   33217 => x"20",
						   33218 => x"34",		-- 0081ec: 3440             MOV.W   #0x2000,R4
						   33219 => x"60",
						   33220 => x"00",		-- 0081ee: 0020            
						   33221 => x"20",
						   33222 => x"36",		-- 0081f0: 3640             MOV.W   #0x2004,R6
						   33223 => x"60",
						   33224 => x"04",		-- 0081f2: 0420            
						   33225 => x"20",
						   33226 => x"A6",		-- 0081f4: A6F4             AND.W   @R4,0x0004(R6)
						   33227 => x"14",
						   33228 => x"04",		-- 0081f6: 0400            
						   33229 => x"00",
						   33230 => x"B0",		-- 0081f8: B0F0             AND.W   #0x2000,Var1
						   33231 => x"10",
						   33232 => x"00",		-- 0081fa: 0020            
						   33233 => x"20",
						   33234 => x"08",		-- 0081fc: 089E            
						   33235 => x"9E",
						   33236 => x"36",		-- 0081fe: 36F5             AND.W   @R5+,R6
						   33237 => x"15",
						   33238 => x"74",		-- 008200: 7440             MOV.B   #0x00aa,R4
						   33239 => x"60",
						   33240 => x"AA",		-- 008202: AA00            
						   33241 => x"00",
						   33242 => x"74",		-- 008204: 74D0             BIS.B   #0x0249,R4
						   33243 => x"F0",
						   33244 => x"49",		-- 008206: 4902            
						   33245 => x"02",
						   33246 => x"05",		-- 008208: 05D4             BIS.W   R4,R5
						   33247 => x"F4",
						   33248 => x"80",		-- 00820a: 80D4             BIS.W   R4,Const2
						   33249 => x"F4",
						   33250 => x"16",		-- 00820c: 169E            
						   33251 => x"9E",
						   33252 => x"15",		-- 00820e: 15D2             BIS.W   &Con1,R5
						   33253 => x"F2",
						   33254 => x"00",		-- 008210: 0020            
						   33255 => x"20",
						   33256 => x"34",		-- 008212: 34D0             BIS.W   #0x2000,R4
						   33257 => x"F0",
						   33258 => x"00",		-- 008214: 0020            
						   33259 => x"20",
						   33260 => x"36",		-- 008216: 36D0             BIS.W   #0x2004,R6
						   33261 => x"F0",
						   33262 => x"04",		-- 008218: 0420            
						   33263 => x"20",
						   33264 => x"A6",		-- 00821a: A6D4             BIS.W   @R4,0x0004(R6)
						   33265 => x"F4",
						   33266 => x"04",		-- 00821c: 0400            
						   33267 => x"00",
						   33268 => x"B0",		-- 00821e: B0D0             BIS.W   #0x2000,Var1
						   33269 => x"F0",
						   33270 => x"00",		-- 008220: 0020            
						   33271 => x"20",
						   33272 => x"E2",		-- 008222: E29D            
						   33273 => x"9D",
						   33274 => x"36",		-- 008224: 36D5             BIS.W   @R5+,R6
						   33275 => x"F5",
						   33276 => x"74",		-- 008226: 7440             MOV.B   #0x00aa,R4
						   33277 => x"60",
						   33278 => x"AA",		-- 008228: AA00            
						   33279 => x"00",
						   33280 => x"74",		-- 00822a: 74E0             XOR.B   #0x0055,R4
						   33281 => x"00",
						   33282 => x"55",		-- 00822c: 5500            
						   33283 => x"00",
						   33284 => x"06",		-- 00822e: 06E5             XOR.W   R5,R6
						   33285 => x"05",
						   33286 => x"80",		-- 008230: 80E4             XOR.W   R4,Const2
						   33287 => x"04",
						   33288 => x"F0",		-- 008232: F09D            
						   33289 => x"9D",
						   33290 => x"15",		-- 008234: 15E2             XOR.W   &Con1,R5
						   33291 => x"02",
						   33292 => x"00",		-- 008236: 0020            
						   33293 => x"20",
						   33294 => x"34",		-- 008238: 3440             MOV.W   #0x2000,R4
						   33295 => x"60",
						   33296 => x"00",		-- 00823a: 0020            
						   33297 => x"20",
						   33298 => x"36",		-- 00823c: 3640             MOV.W   #0x2004,R6
						   33299 => x"60",
						   33300 => x"04",		-- 00823e: 0420            
						   33301 => x"20",
						   33302 => x"A6",		-- 008240: A6E4             XOR.W   @R4,0x0004(R6)
						   33303 => x"04",
						   33304 => x"04",		-- 008242: 0400            
						   33305 => x"00",
						   33306 => x"B0",		-- 008244: B0E0             XOR.W   #0x2000,Var1
						   33307 => x"00",
						   33308 => x"00",		-- 008246: 0020            
						   33309 => x"20",
						   33310 => x"BC",		-- 008248: BC9D            
						   33311 => x"9D",
						   33312 => x"36",		-- 00824a: 36E5             XOR.W   @R5+,R6
						   33313 => x"05",
						   33314 => x"74",		-- 00824c: 7440             MOV.B   #0x00aa,R4
						   33315 => x"60",
						   33316 => x"AA",		-- 00824e: AA00            
						   33317 => x"00",
						   33318 => x"74",		-- 008250: 74D0             BIS.B   #0x0249,R4
						   33319 => x"F0",
						   33320 => x"49",		-- 008252: 4902            
						   33321 => x"02",
						   33322 => x"05",		-- 008254: 05D4             BIS.W   R4,R5
						   33323 => x"F4",
						   33324 => x"80",		-- 008256: 80D4             BIS.W   R4,Const2
						   33325 => x"F4",
						   33326 => x"CA",		-- 008258: CA9D            
						   33327 => x"9D",
						   33328 => x"15",		-- 00825a: 15D2             BIS.W   &Con1,R5
						   33329 => x"F2",
						   33330 => x"00",		-- 00825c: 0020            
						   33331 => x"20",
						   33332 => x"34",		-- 00825e: 3440             MOV.W   #0x2000,R4
						   33333 => x"60",
						   33334 => x"00",		-- 008260: 0020            
						   33335 => x"20",
						   33336 => x"36",		-- 008262: 3640             MOV.W   #0x2004,R6
						   33337 => x"60",
						   33338 => x"04",		-- 008264: 0420            
						   33339 => x"20",
						   33340 => x"A6",		-- 008266: A6D4             BIS.W   @R4,0x0004(R6)
						   33341 => x"F4",
						   33342 => x"04",		-- 008268: 0400            
						   33343 => x"00",
						   33344 => x"B0",		-- 00826a: B0D0             BIS.W   #0x2000,Var1
						   33345 => x"F0",
						   33346 => x"00",		-- 00826c: 0020            
						   33347 => x"20",
						   33348 => x"96",		-- 00826e: 969D            
						   33349 => x"9D",
						   33350 => x"36",		-- 008270: 36D5             BIS.W   @R5+,R6
						   33351 => x"F5",
						   33352 => x"74",		-- 008272: 7440             MOV.B   #0x00aa,R4
						   33353 => x"60",
						   33354 => x"AA",		-- 008274: AA00            
						   33355 => x"00",
						   33356 => x"74",		-- 008276: 74C0             BIC.B   #0x0018,R4
						   33357 => x"E0",
						   33358 => x"18",		-- 008278: 1800            
						   33359 => x"00",
						   33360 => x"05",		-- 00827a: 05C4             BIC.W   R4,R5
						   33361 => x"E4",
						   33362 => x"80",		-- 00827c: 80C4             BIC.W   R4,Const2
						   33363 => x"E4",
						   33364 => x"A4",		-- 00827e: A49D            
						   33365 => x"9D",
						   33366 => x"15",		-- 008280: 15C2             BIC.W   &Con1,R5
						   33367 => x"E2",
						   33368 => x"00",		-- 008282: 0020            
						   33369 => x"20",
						   33370 => x"34",		-- 008284: 3440             MOV.W   #0x2000,R4
						   33371 => x"60",
						   33372 => x"00",		-- 008286: 0020            
						   33373 => x"20",
						   33374 => x"36",		-- 008288: 3640             MOV.W   #0x2004,R6
						   33375 => x"60",
						   33376 => x"04",		-- 00828a: 0420            
						   33377 => x"20",
						   33378 => x"A6",		-- 00828c: A6C4             BIC.W   @R4,0x0004(R6)
						   33379 => x"E4",
						   33380 => x"04",		-- 00828e: 0400            
						   33381 => x"00",
						   33382 => x"B0",		-- 008290: B0C0             BIC.W   #0x2000,Var1
						   33383 => x"E0",
						   33384 => x"00",		-- 008292: 0020            
						   33385 => x"20",
						   33386 => x"70",		-- 008294: 709D            
						   33387 => x"9D",
						   33388 => x"36",		-- 008296: 36C5             BIC.W   @R5+,R6
						   33389 => x"E5",
						   33390 => x"74",		-- 008298: 7440             MOV.B   #0x00aa,R4
						   33391 => x"60",
						   33392 => x"AA",		-- 00829a: AA00            
						   33393 => x"00",
						   33394 => x"74",		-- 00829c: 74B0             BIT.B   #0x0018,R4
						   33395 => x"D0",
						   33396 => x"18",		-- 00829e: 1800            
						   33397 => x"00",
						   33398 => x"05",		-- 0082a0: 05B4             BIT.W   R4,R5
						   33399 => x"D4",
						   33400 => x"80",		-- 0082a2: 80B4             BIT.W   R4,Const2
						   33401 => x"D4",
						   33402 => x"7E",		-- 0082a4: 7E9D            
						   33403 => x"9D",
						   33404 => x"15",		-- 0082a6: 15B2             BIT.W   &Con1,R5
						   33405 => x"D2",
						   33406 => x"00",		-- 0082a8: 0020            
						   33407 => x"20",
						   33408 => x"34",		-- 0082aa: 3440             MOV.W   #0x2000,R4
						   33409 => x"60",
						   33410 => x"00",		-- 0082ac: 0020            
						   33411 => x"20",
						   33412 => x"36",		-- 0082ae: 3640             MOV.W   #0x2004,R6
						   33413 => x"60",
						   33414 => x"04",		-- 0082b0: 0420            
						   33415 => x"20",
						   33416 => x"A6",		-- 0082b2: A6B4             BIT.W   @R4,0x0004(R6)
						   33417 => x"D4",
						   33418 => x"04",		-- 0082b4: 0400            
						   33419 => x"00",
						   33420 => x"B0",		-- 0082b6: B0B0             BIT.W   #0x2000,Var1
						   33421 => x"D0",
						   33422 => x"00",		-- 0082b8: 0020            
						   33423 => x"20",
						   33424 => x"4A",		-- 0082ba: 4A9D            
						   33425 => x"9D",
						   33426 => x"36",		-- 0082bc: 36B5             BIT.W   @R5+,R6
						   33427 => x"D5",
						   33428 => x"75",		-- 0082be: 7540             MOV.B   #0x0063,R5
						   33429 => x"60",
						   33430 => x"63",		-- 0082c0: 6300            
						   33431 => x"00",
						   33432 => x"75",		-- 0082c2: 7590             CMP.B   #0x0063,R5
						   33433 => x"B0",
						   33434 => x"63",		-- 0082c4: 6300            
						   33435 => x"00",
						   33436 => x"75",		-- 0082c6: 7590             CMP.B   #0x004d,R5
						   33437 => x"B0",
						   33438 => x"4D",		-- 0082c8: 4D00            
						   33439 => x"00",
						   33440 => x"05",		-- 0082ca: 0594             CMP.W   R4,R5
						   33441 => x"B4",
						   33442 => x"80",		-- 0082cc: 8094             CMP.W   R4,Const2
						   33443 => x"B4",
						   33444 => x"54",		-- 0082ce: 549D            
						   33445 => x"9D",
						   33446 => x"15",		-- 0082d0: 1592             CMP.W   &Con1,R5
						   33447 => x"B2",
						   33448 => x"00",		-- 0082d2: 0020            
						   33449 => x"20",
						   33450 => x"34",		-- 0082d4: 3440             MOV.W   #0x2000,R4
						   33451 => x"60",
						   33452 => x"00",		-- 0082d6: 0020            
						   33453 => x"20",
						   33454 => x"36",		-- 0082d8: 3640             MOV.W   #0x2004,R6
						   33455 => x"60",
						   33456 => x"04",		-- 0082da: 0420            
						   33457 => x"20",
						   33458 => x"A6",		-- 0082dc: A694             CMP.W   @R4,0x0004(R6)
						   33459 => x"B4",
						   33460 => x"04",		-- 0082de: 0400            
						   33461 => x"00",
						   33462 => x"B0",		-- 0082e0: B090             CMP.W   #0x2000,Var1
						   33463 => x"B0",
						   33464 => x"00",		-- 0082e2: 0020            
						   33465 => x"20",
						   33466 => x"20",		-- 0082e4: 209D            
						   33467 => x"9D",
						   33468 => x"36",		-- 0082e6: 3695             CMP.W   @R5+,R6
						   33469 => x"B5",
						   33470 => x"77",		-- 0082e8: 7740             MOV.B   #0xff9d,R7
						   33471 => x"60",
						   33472 => x"9D",		-- 0082ea: 9DFF            
						   33473 => x"FF",
						   33474 => x"04",		-- 0082f2: 0493             TST.W   R4
						   33475 => x"B3",
						   33476 => x"80",		-- 0082f4: 8093             TST.W   Const2
						   33477 => x"B3",
						   33478 => x"2C",		-- 0082f6: 2C9D            
						   33479 => x"9D",
						   33480 => x"82",		-- 0082f8: 8293             TST.W   &Con1
						   33481 => x"B3",
						   33482 => x"00",		-- 0082fa: 0020            
						   33483 => x"20",
						   33484 => x"B0",		-- 0082fc: B040             MOV.W   #0x2000,Var1
						   33485 => x"60",
						   33486 => x"00",		-- 0082fe: 0020            
						   33487 => x"20",
						   33488 => x"04",		-- 008300: 049D            
						   33489 => x"9D",
						   33490 => x"34",		-- 008302: 3440             MOV.W   #0x2000,R4
						   33491 => x"60",
						   33492 => x"00",		-- 008304: 0020            
						   33493 => x"20",
						   33494 => x"80",		-- 008306: 8093             TST.W   Var1
						   33495 => x"B3",
						   33496 => x"FC",		-- 008308: FC9C            
						   33497 => x"9C",
						   33498 => x"84",		-- 00830a: 8493             TST.W   0x0004(R4)
						   33499 => x"B3",
						   33500 => x"04",		-- 00830c: 0400            
						   33501 => x"00",
						   33502 => x"54",		-- 00830e: 5443             MOV.B   #1,R4
						   33503 => x"63",
						   33504 => x"90",		-- 008316: 9050             ADD.W   Const2,Const2
						   33505 => x"70",
						   33506 => x"0A",		-- 008318: 0A9D            
						   33507 => x"9D",
						   33508 => x"08",		-- 00831a: 089D            
						   33509 => x"9D",
						   33510 => x"00",		-- 00831e: 0020            
						   33511 => x"20",
						   33512 => x"00",		-- 008320: 0020            
						   33513 => x"20",
						   33514 => x"B0",		-- 008322: B040             MOV.W   #0x2000,Var1
						   33515 => x"60",
						   33516 => x"00",		-- 008324: 0020            
						   33517 => x"20",
						   33518 => x"DE",		-- 008326: DE9C            
						   33519 => x"9C",
						   33520 => x"34",		-- 008328: 3440             MOV.W   #0x2000,R4
						   33521 => x"60",
						   33522 => x"00",		-- 00832a: 0020            
						   33523 => x"20",
						   33524 => x"90",		-- 00832c: 9050             ADD.W   Var1,Var1
						   33525 => x"70",
						   33526 => x"D6",		-- 00832e: D69C            
						   33527 => x"9C",
						   33528 => x"D4",		-- 008330: D49C            
						   33529 => x"9C",
						   33530 => x"04",		-- 008334: 0400            
						   33531 => x"00",
						   33532 => x"04",		-- 008336: 0400            
						   33533 => x"00",
						   33534 => x"74",		-- 008338: 7440             MOV.B   #0x0020,R4
						   33535 => x"60",
						   33536 => x"20",		-- 00833a: 2000            
						   33537 => x"00",
						   33538 => x"44",		-- 00833c: 4411             RRA.B   R4
						   33539 => x"31",
						   33540 => x"44",		-- 00833e: 4411             RRA.B   R4
						   33541 => x"31",
						   33542 => x"DE",		-- 008344: DE9C            
						   33543 => x"9C",
						   33544 => x"00",		-- 008348: 0020            
						   33545 => x"20",
						   33546 => x"B0",		-- 00834a: B040             MOV.W   #0x2000,Var1
						   33547 => x"60",
						   33548 => x"00",		-- 00834c: 0020            
						   33549 => x"20",
						   33550 => x"B6",		-- 00834e: B69C            
						   33551 => x"9C",
						   33552 => x"34",		-- 008350: 3440             MOV.W   #0x2000,R4
						   33553 => x"60",
						   33554 => x"00",		-- 008352: 0020            
						   33555 => x"20",
						   33556 => x"AE",		-- 008356: AE9C            
						   33557 => x"9C",
						   33558 => x"04",		-- 00835a: 0400            
						   33559 => x"00",
						   33560 => x"77",		-- 00835e: 7740             MOV.B   #0x0080,R7
						   33561 => x"60",
						   33562 => x"80",		-- 008360: 8000            
						   33563 => x"00",
						   33564 => x"90",		-- 008368: 9060             ADDC.W  Const2,Const2
						   33565 => x"80",
						   33566 => x"B8",		-- 00836a: B89C            
						   33567 => x"9C",
						   33568 => x"B6",		-- 00836c: B69C            
						   33569 => x"9C",
						   33570 => x"00",		-- 008370: 0020            
						   33571 => x"20",
						   33572 => x"00",		-- 008372: 0020            
						   33573 => x"20",
						   33574 => x"B0",		-- 008374: B040             MOV.W   #0x2000,Var1
						   33575 => x"60",
						   33576 => x"00",		-- 008376: 0020            
						   33577 => x"20",
						   33578 => x"8C",		-- 008378: 8C9C            
						   33579 => x"9C",
						   33580 => x"34",		-- 00837a: 3440             MOV.W   #0x2000,R4
						   33581 => x"60",
						   33582 => x"00",		-- 00837c: 0020            
						   33583 => x"20",
						   33584 => x"90",		-- 00837e: 9060             ADDC.W  Var1,Var1
						   33585 => x"80",
						   33586 => x"84",		-- 008380: 849C            
						   33587 => x"9C",
						   33588 => x"82",		-- 008382: 829C            
						   33589 => x"9C",
						   33590 => x"04",		-- 008386: 0400            
						   33591 => x"00",
						   33592 => x"04",		-- 008388: 0400            
						   33593 => x"00",
						   33594 => x"58",		-- 00838c: 5843             MOV.B   #1,R8
						   33595 => x"63",
						   33596 => x"48",		-- 00838e: 4810             RRC.B   R8
						   33597 => x"30",
						   33598 => x"48",		-- 008390: 4810             RRC.B   R8
						   33599 => x"30",
						   33600 => x"8C",		-- 008396: 8C9C            
						   33601 => x"9C",
						   33602 => x"00",		-- 00839a: 0020            
						   33603 => x"20",
						   33604 => x"B0",		-- 00839c: B040             MOV.W   #0x2000,Var1
						   33605 => x"60",
						   33606 => x"00",		-- 00839e: 0020            
						   33607 => x"20",
						   33608 => x"64",		-- 0083a0: 649C            
						   33609 => x"9C",
						   33610 => x"34",		-- 0083a2: 3440             MOV.W   #0x2000,R4
						   33611 => x"60",
						   33612 => x"00",		-- 0083a4: 0020            
						   33613 => x"20",
						   33614 => x"5C",		-- 0083a8: 5C9C            
						   33615 => x"9C",
						   33616 => x"04",		-- 0083ac: 0400            
						   33617 => x"00",
						   33618 => x"34",		-- 0083ae: 3440             MOV.W   #0x00ff,R4
						   33619 => x"60",
						   33620 => x"FF",		-- 0083b0: FF00            
						   33621 => x"00",
						   33622 => x"6C",		-- 0083b6: 6C9C            
						   33623 => x"9C",
						   33624 => x"00",		-- 0083ba: 0020            
						   33625 => x"20",
						   33626 => x"B0",		-- 0083bc: B040             MOV.W   #0x2000,Var1
						   33627 => x"60",
						   33628 => x"00",		-- 0083be: 0020            
						   33629 => x"20",
						   33630 => x"44",		-- 0083c0: 449C            
						   33631 => x"9C",
						   33632 => x"34",		-- 0083c2: 3440             MOV.W   #0x2000,R4
						   33633 => x"60",
						   33634 => x"00",		-- 0083c4: 0020            
						   33635 => x"20",
						   33636 => x"3C",		-- 0083c8: 3C9C            
						   33637 => x"9C",
						   33638 => x"04",		-- 0083cc: 0400            
						   33639 => x"00",
						   33640 => x"34",		-- 0083ce: 3440             MOV.W   #0x00ff,R4
						   33641 => x"60",
						   33642 => x"FF",		-- 0083d0: FF00            
						   33643 => x"00",
						   33644 => x"4C",		-- 0083d6: 4C9C            
						   33645 => x"9C",
						   33646 => x"00",		-- 0083da: 0020            
						   33647 => x"20",
						   33648 => x"B0",		-- 0083dc: B040             MOV.W   #0x2000,Var1
						   33649 => x"60",
						   33650 => x"00",		-- 0083de: 0020            
						   33651 => x"20",
						   33652 => x"24",		-- 0083e0: 249C            
						   33653 => x"9C",
						   33654 => x"34",		-- 0083e2: 3440             MOV.W   #0x2000,R4
						   33655 => x"60",
						   33656 => x"00",		-- 0083e4: 0020            
						   33657 => x"20",
						   33658 => x"1C",		-- 0083e8: 1C9C            
						   33659 => x"9C",
						   33660 => x"04",		-- 0083ec: 0400            
						   33661 => x"00",
						   33662 => x"3A",		-- 0083fa: 3A40             MOV.W   #0x001c,R10
						   33663 => x"60",
						   33664 => x"1C",		-- 0083fc: 1C00            
						   33665 => x"00",
						   33666 => x"0A",		-- 0083fe: 0A43             CLR.W   R10
						   33667 => x"63",
						   33668 => x"80",		-- 008400: 8043             CLR.W   Var1
						   33669 => x"63",
						   33670 => x"02",		-- 008402: 029C            
						   33671 => x"9C",
						   33672 => x"82",		-- 008404: 8243             CLR.W   &Con1
						   33673 => x"63",
						   33674 => x"00",		-- 008406: 0020            
						   33675 => x"20",
						   33676 => x"3A",		-- 008408: 3A40             MOV.W   #0x2000,R10
						   33677 => x"60",
						   33678 => x"00",		-- 00840a: 0020            
						   33679 => x"20",
						   33680 => x"8A",		-- 00840c: 8A43             CLR.W   0x0002(R10)
						   33681 => x"63",
						   33682 => x"02",		-- 00840e: 0200            
						   33683 => x"00",
						   33684 => x"00",		-- 008422: 0024             JEQ     (_jeq)
						   33685 => x"44",
						   33686 => x"FE",		-- 008426: FE27             JEQ     (_jeq)
						   33687 => x"47",
						   33688 => x"00",		-- 00842a: 0024             JEQ     (_jz)
						   33689 => x"44",
						   33690 => x"FE",		-- 00842e: FE27             JEQ     (_jz)
						   33691 => x"47",
						   33692 => x"14",		-- 008430: 1443             MOV.W   #1,R4
						   33693 => x"63",
						   33694 => x"04",		-- 008432: 0493             TST.W   R4
						   33695 => x"B3",
						   33696 => x"00",		-- 008434: 0034             JGE     (_jge)
						   33697 => x"54",
						   33698 => x"04",		-- 008436: 0443             CLR.W   R4
						   33699 => x"63",
						   33700 => x"14",		-- 008438: 1493             CMP.W   #1,R4
						   33701 => x"B3",
						   33702 => x"FD",		-- 00843a: FD37             JGE     (_jge)
						   33703 => x"57",
						   33704 => x"04",		-- 00843c: 0443             CLR.W   R4
						   33705 => x"63",
						   33706 => x"14",		-- 00843e: 1493             CMP.W   #1,R4
						   33707 => x"B3",
						   33708 => x"00",		-- 008440: 0038             JL      (_jl)
						   33709 => x"58",
						   33710 => x"14",		-- 008442: 1443             MOV.W   #1,R4
						   33711 => x"63",
						   33712 => x"04",		-- 008444: 0493             TST.W   R4
						   33713 => x"B3",
						   33714 => x"FD",		-- 008446: FD3B             JL      (_jl)
						   33715 => x"5B",
						   33716 => x"00",		-- 008448: 003C             JMP     (_jmp)
						   33717 => x"5C",
						   33718 => x"03",		-- 00844a: 0343             NOP     
						   33719 => x"63",
						   33720 => x"00",		-- 00844e: 0030             JN      (_jn)
						   33721 => x"50",
						   33722 => x"FE",		-- 008452: FE33             JN      (_jn)
						   33723 => x"53",
						   33724 => x"00",		-- 008466: 0020             JNE     (_jne)
						   33725 => x"40",
						   33726 => x"FE",		-- 00846a: FE23             JNE     (_jne)
						   33727 => x"43",
						   33728 => x"00",		-- 00846e: 0020             JNE     (_jnz)
						   33729 => x"40",
						   33730 => x"FE",		-- 008472: FE23             JNE     (_jnz)
						   33731 => x"43",
						   33732 => x"34",		-- 008474: 3440             MOV.W   #0x847a,R4
						   33733 => x"60",
						   33734 => x"7A",		-- 008476: 7A84            
						   33735 => x"84",
						   33736 => x"B0",		-- 00847a: B040             MOV.W   #0x8484,Const2
						   33737 => x"60",
						   33738 => x"84",		-- 00847c: 8484            
						   33739 => x"84",
						   33740 => x"A4",		-- 00847e: A49B            
						   33741 => x"9B",
						   33742 => x"A0",		-- 008482: A09B            
						   33743 => x"9B",
						   33744 => x"88",		-- 008486: 8884            
						   33745 => x"84",
						   33746 => x"03",		-- 008488: 0343             NOP     
						   33747 => x"63",
						   33748 => x"34",		-- 00848a: 3440             MOV.W   #0x00ff,R4
						   33749 => x"60",
						   33750 => x"FF",		-- 00848c: FF00            
						   33751 => x"00",
						   33752 => x"F0",		-- 008490: F0F0            
						   33753 => x"F0",
						   33754 => x"00",		-- 008496: 0020            
						   33755 => x"20",
						   33756 => x"34",		-- 008498: 3440             MOV.W   #0x2000,R4
						   33757 => x"60",
						   33758 => x"00",		-- 00849a: 0020            
						   33759 => x"20",
						   33760 => x"00",		-- 00849e: 0000            
						   33761 => x"00",
						   33762 => x"00",		-- 0084a2: 0020            
						   33763 => x"20",
						   33764 => x"78",		-- 0084aa: 789B            
						   33765 => x"9B",
						   33766 => x"00",		-- 0084ae: 0020            
						   33767 => x"20",
						   33768 => x"B0",		-- 0084b0: B040             MOV.W   #0x2000,Var1
						   33769 => x"60",
						   33770 => x"00",		-- 0084b2: 0020            
						   33771 => x"20",
						   33772 => x"50",		-- 0084b4: 509B            
						   33773 => x"9B",
						   33774 => x"34",		-- 0084b6: 3440             MOV.W   #0x2000,R4
						   33775 => x"60",
						   33776 => x"00",		-- 0084b8: 0020            
						   33777 => x"20",
						   33778 => x"48",		-- 0084bc: 489B            
						   33779 => x"9B",
						   33780 => x"04",		-- 0084c0: 0400            
						   33781 => x"00",
						   33782 => x"05",		-- 0084c4: 0543             CLR.W   R5
						   33783 => x"63",
						   33784 => x"34",		-- 0084c6: 3440             MOV.W   #0x84e4,R4
						   33785 => x"60",
						   33786 => x"E4",		-- 0084c8: E484            
						   33787 => x"84",
						   33788 => x"B0",		-- 0084ca: B040             MOV.W   #0x84e4,Var1
						   33789 => x"60",
						   33790 => x"E4",		-- 0084cc: E484            
						   33791 => x"84",
						   33792 => x"36",		-- 0084ce: 369B            
						   33793 => x"9B",
						   33794 => x"E4",		-- 0084d2: E484            
						   33795 => x"84",
						   33796 => x"2C",		-- 0084d8: 2C9B            
						   33797 => x"9B",
						   33798 => x"E4",		-- 0084dc: E484            
						   33799 => x"84",
						   33800 => x"3E",		-- 0084e0: 3E80            
						   33801 => x"80",
						   33802 => x"03",		-- 0084e2: 0343             NOP     
						   33803 => x"63",
						   33804 => x"35",		-- 0084e4: 3550             ADD.W   #0x0003,R5
						   33805 => x"70",
						   33806 => x"03",		-- 0084e6: 0300            
						   33807 => x"00",
						   33808 => x"F2",		-- 0084ea: F2E0             XOR.B   #0x0040,&P6OUT
						   33809 => x"00",
						   33810 => x"40",		-- 0084ec: 4000            
						   33811 => x"00",
						   33812 => x"43",		-- 0084ee: 4302            
						   33813 => x"02",
						   33814 => x"E2",		-- 0084f0: E2C3             BIC.B   #2,&P4IFG
						   33815 => x"E3",
						   33816 => x"3D",		-- 0084f2: 3D02            
						   33817 => x"02",
						   33818 => x"32",		-- 0084f6: 32D0             BIS.W   #0x0010,SR
						   33819 => x"F0",
        -- IRQ Vectors (Interrupts)
                           65534 =>  x"00",		-- Reset Vector = xFFFE:xFFFF
                           65535 =>  x"80",		--  Startup Value = x8000

                           others => x"00");

    signal EN : std_logic;

    begin
    -- Note 1:  The bus system uses a 16-bit Address (MAB)
    --          This address size can access locations from x0000 to xFFFF
    --          But our array is only defined from x8000 to xFFFF and
    --          if we try to access it with any other address, it will crash.
    --          So the first thing we need to do is create a local enable that
    --          will only assert when MAB is within x8000 to xFFFF.

     LOCAL_EN : process (MAB) 
       begin
         if ( (to_integer(unsigned(MAB)) >= 32768) and (to_integer(unsigned(MAB)) <= 65535)) then
           EN <= '1';
         else 
           EN <= '0';
        end if;
      end process;


    -- Note 2:  The bus system uses a 16-bit Address (MAB)
    --          The MDB_out is also provided as a 16-bit word
    --          However, the memory array is actually built as 8-bit bytes.
    --          So for a given 16-bit MAB, we give MDB_out = HB : LB
    --                                                 or  = ROM(MAB);1) : ROM(MAB)

    MEMORY_ROM : process (clk) 
     begin
        if (rising_edge(clk)) then
            if (EN='1' and write='0') then                      
              MDB_in <= ROM(to_integer(unsigned(MAB)) + 1 ) & ROM(to_integer(unsigned(MAB))); 
            end if;
      end if;
   end process;


end architecture;