library IEEE;
    use IEEE.std_logic_1164.all;
    use IEEE.numeric_std.all;
    package lowlife is
    constant FORMAT_2 : integer := 1;
    constant JMP1 : integer := 2;
    constant JMP2 : integer := 3;
    constant MOV : integer := 4;
    constant OFFSET : integer := 0;
    end lowlife;
