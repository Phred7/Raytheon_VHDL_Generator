library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;


entity baseline_memory is
    port ( clk	: in	std_logic;
         MAB		: in	std_logic_vector(15 downto 0);
         MDB_in  	: out	std_logic_vector(15 downto 0);
         MDB_out  	: in	std_logic_vector(15 downto 0);
         write	    : in	std_logic);
end entity;

architecture baseline_memory_arch of baseline_memory is

type rom_type is array (32768 to 65535) of std_logic_vector(7 downto 0);  -- this is MAB: x8000 to xFFFF
    
constant ROM : rom_type :=(						   50246 => x"B2",		-- 00c446: B240             MOV.W   #0x5a80,&WDTCTL_L
						   50247 => x"40",
						   50248 => x"80",		-- 00c448: 805A            
						   50249 => x"5A",
						   50250 => x"CC",		-- 00c44a: CC01            
						   50251 => x"01",
						   50252 => x"91",		-- 00c44c: 9142             MOV.W   &$P$T0$1,0x0002(SP)
						   50253 => x"42",
						   50254 => x"5C",		-- 00c44e: 5C86            
						   50255 => x"86",
						   50256 => x"02",		-- 00c450: 0200            
						   50257 => x"00",
						   50258 => x"91",		-- 00c452: 9142             MOV.W   &0x865e,0x0004(SP)
						   50259 => x"42",
						   50260 => x"5E",		-- 00c454: 5E86            
						   50261 => x"86",
						   50262 => x"04",		-- 00c456: 0400            
						   50263 => x"00",
						   50264 => x"91",		-- 00c458: 9142             MOV.W   &0x8660,0x0006(SP)
						   50265 => x"42",
						   50266 => x"60",		-- 00c45a: 6086            
						   50267 => x"86",
						   50268 => x"06",		-- 00c45c: 0600            
						   50269 => x"00",
						   50270 => x"91",		-- 00c45e: 9142             MOV.W   &0x8662,0x0008(SP)
						   50271 => x"42",
						   50272 => x"62",		-- 00c460: 6286            
						   50273 => x"86",
						   50274 => x"08",		-- 00c462: 0800            
						   50275 => x"00",
						   50276 => x"81",		-- 00c464: 8143             CLR.W   0x000c(SP)
						   50277 => x"43",
						   50278 => x"0C",		-- 00c466: 0C00            
						   50279 => x"00",
						   50280 => x"1C",		-- 00c468: 1C41             MOV.W   0x000a(SP),R12
						   50281 => x"41",
						   50282 => x"0A",		-- 00c46a: 0A00            
						   50283 => x"00",
						   50284 => x"B0",		-- 00c46c: B012             CALL    #buff_value
						   50285 => x"12",
						   50286 => x"54",		-- 00c46e: 54CD            
						   50287 => x"CD",
						   50288 => x"1C",		-- 00c470: 1C41             MOV.W   0x000e(SP),R12
						   50289 => x"41",
						   50290 => x"0E",		-- 00c472: 0E00            
						   50291 => x"00",
						   50292 => x"B0",		-- 00c474: B012             CALL    #buff_value
						   50293 => x"12",
						   50294 => x"54",		-- 00c476: 54CD            
						   50295 => x"CD",
						   50296 => x"81",		-- 00c478: 8193             TST.W   0x000c(SP)
						   50297 => x"93",
						   50298 => x"0C",		-- 00c47a: 0C00            
						   50299 => x"00",
						   50300 => x"07",		-- 00c47c: 0720             JNE     ($C$L1)
						   50301 => x"20",
						   50302 => x"0F",		-- 00c47e: 0F41             MOV.W   SP,R15
						   50303 => x"41",
						   50304 => x"2F",		-- 00c480: 2F53             INCD.W  R15
						   50305 => x"53",
						   50306 => x"81",		-- 00c482: 814F             MOV.W   R15,0x0000(SP)
						   50307 => x"4F",
						   50308 => x"00",		-- 00c484: 0000            
						   50309 => x"00",
						   50310 => x"B0",		-- 00c486: B012             CALL    #printf
						   50311 => x"12",
						   50312 => x"1E",		-- 00c488: 1EC9            
						   50313 => x"C9",
						   50314 => x"05",		-- 00c48a: 053C             JMP     ($C$L2)
						   50315 => x"3C",
						   50316 => x"B1",		-- 00c48c: B140             MOV.W   #0x8654,0x0000(SP)
						   50317 => x"40",
						   50318 => x"54",		-- 00c48e: 5486            
						   50319 => x"86",
						   50320 => x"00",		-- 00c490: 0000            
						   50321 => x"00",
						   50322 => x"B0",		-- 00c492: B012             CALL    #printf
						   50323 => x"12",
						   50324 => x"1E",		-- 00c494: 1EC9            
						   50325 => x"C9",
						   50326 => x"0C",		-- 00c496: 0C43             CLR.W   R12
						   50327 => x"43",
						   50328 => x"31",		-- 00c498: 3150             ADD.W   #0x0010,SP
						   50329 => x"50",
						   50330 => x"10",		-- 00c49a: 1000            
						   50331 => x"00",
						   50332 => x"30",		-- 00c49c: 3041             RET     
						   50333 => x"41",
						   -- Begin: getdevice
						   50334 => x"0A",		-- 00c49e: 0A12             PUSH    R10
						   50335 => x"12",
						   50336 => x"09",		-- 00c4a0: 0912             PUSH    R9
						   50337 => x"12",
						   50338 => x"08",		-- 00c4a2: 0812             PUSH    R8
						   50339 => x"12",
						   50340 => x"31",		-- 00c4a4: 3180             SUB.W   #0x000a,SP
						   50341 => x"80",
						   50342 => x"0A",		-- 00c4a6: 0A00            
						   50343 => x"00",
						   50344 => x"08",		-- 00c4a8: 084C             MOV.W   R12,R8
						   50345 => x"4C",
						   50346 => x"2C",		-- 00c4aa: 2C48             MOV.W   @R8,R12
						   50347 => x"48",
						   50348 => x"3D",		-- 00c4ac: 3D40             MOV.W   #0x003a,R13
						   50349 => x"40",
						   50350 => x"3A",		-- 00c4ae: 3A00            
						   50351 => x"00",
						   50352 => x"B0",		-- 00c4b0: B012             CALL    #strchr
						   50353 => x"12",
						   50354 => x"A8",		-- 00c4b2: A8CC            
						   50355 => x"CC",
						   50356 => x"09",		-- 00c4b4: 094C             MOV.W   R12,R9
						   50357 => x"4C",
						   50358 => x"09",		-- 00c4b6: 0993             TST.W   R9
						   50359 => x"93",
						   50360 => x"18",		-- 00c4b8: 1824             JEQ     ($C$L5)
						   50361 => x"24",
						   50362 => x"0A",		-- 00c4ba: 0A49             MOV.W   R9,R10
						   50363 => x"49",
						   50364 => x"2A",		-- 00c4bc: 2A88             SUB.W   @R8,R10
						   50365 => x"88",
						   50366 => x"3A",		-- 00c4be: 3A90             CMP.W   #0x0009,R10
						   50367 => x"90",
						   50368 => x"09",		-- 00c4c0: 0900            
						   50369 => x"00",
						   50370 => x"01",		-- 00c4c2: 0138             JL      ($C$L4)
						   50371 => x"38",
						   50372 => x"3A",		-- 00c4c4: 3A42             MOV.W   #8,R10
						   50373 => x"42",
						   50374 => x"2D",		-- 00c4c6: 2D48             MOV.W   @R8,R13
						   50375 => x"48",
						   50376 => x"0E",		-- 00c4c8: 0E4A             MOV.W   R10,R14
						   50377 => x"4A",
						   50378 => x"0C",		-- 00c4ca: 0C41             MOV.W   SP,R12
						   50379 => x"41",
						   50380 => x"B0",		-- 00c4cc: B012             CALL    #strncpy
						   50381 => x"12",
						   50382 => x"D0",		-- 00c4ce: D0CA            
						   50383 => x"CA",
						   50384 => x"0F",		-- 00c4d0: 0F41             MOV.W   SP,R15
						   50385 => x"41",
						   50386 => x"0F",		-- 00c4d2: 0F5A             ADD.W   R10,R15
						   50387 => x"5A",
						   50388 => x"CF",		-- 00c4d4: CF43             CLR.B   0x0000(R15)
						   50389 => x"43",
						   50390 => x"00",		-- 00c4d6: 0000            
						   50391 => x"00",
						   50392 => x"0C",		-- 00c4d8: 0C41             MOV.W   SP,R12
						   50393 => x"41",
						   50394 => x"B0",		-- 00c4da: B012             CALL    #finddevice
						   50395 => x"12",
						   50396 => x"8E",		-- 00c4dc: 8EC9            
						   50397 => x"C9",
						   50398 => x"0C",		-- 00c4de: 0C93             TST.W   R12
						   50399 => x"93",
						   50400 => x"04",		-- 00c4e0: 0424             JEQ     ($C$L5)
						   50401 => x"24",
						   50402 => x"19",		-- 00c4e2: 1953             INC.W   R9
						   50403 => x"53",
						   50404 => x"88",		-- 00c4e4: 8849             MOV.W   R9,0x0000(R8)
						   50405 => x"49",
						   50406 => x"00",		-- 00c4e6: 0000            
						   50407 => x"00",
						   50408 => x"02",		-- 00c4e8: 023C             JMP     ($C$L6)
						   50409 => x"3C",
						   50410 => x"3C",		-- 00c4ea: 3C40             MOV.W   #0x2078,R12
						   50411 => x"40",
						   50412 => x"78",		-- 00c4ec: 7820            
						   50413 => x"20",
						   50414 => x"31",		-- 00c4ee: 3150             ADD.W   #0x000a,SP
						   50415 => x"50",
						   50416 => x"0A",		-- 00c4f0: 0A00            
						   50417 => x"00",
						   50418 => x"30",		-- 00c4f2: 3040             BR      #__mspabi_func_epilog_3
						   50419 => x"40",
						   50420 => x"A4",		-- 00c4f4: A4CD            
						   50421 => x"CD",
						   -- Begin: __mspabi_divul
						   -- Begin: __mspabi_remul
						   50422 => x"0A",		-- 00c4f6: 0A12             PUSH    R10
						   50423 => x"12",
						   50424 => x"09",		-- 00c4f8: 0912             PUSH    R9
						   50425 => x"12",
						   50426 => x"09",		-- 00c4fa: 0943             CLR.W   R9
						   50427 => x"43",
						   50428 => x"0A",		-- 00c4fc: 0A43             CLR.W   R10
						   50429 => x"43",
						   50430 => x"1B",		-- 00c4fe: 1B43             MOV.W   #1,R11
						   50431 => x"43",
						   50432 => x"0F",		-- 00c500: 0F93             TST.W   R15
						   50433 => x"93",
						   50434 => x"04",		-- 00c502: 0424             JEQ     (div_loop_lo)
						   50435 => x"24",
						   50436 => x"09",		-- 00c504: 094D             MOV.W   R13,R9
						   50437 => x"4D",
						   50438 => x"0D",		-- 00c506: 0D4C             MOV.W   R12,R13
						   50439 => x"4C",
						   50440 => x"0C",		-- 00c508: 0C43             CLR.W   R12
						   50441 => x"43",
						   50442 => x"0D",		-- 00c50a: 0D3C             JMP     (div_loop_hi)
						   50443 => x"3C",
						   -- Begin: div_loop_lo
						   50444 => x"0C",		-- 00c50c: 0C5C             RLA.W   R12
						   50445 => x"5C",
						   50446 => x"0D",		-- 00c50e: 0D6D             RLC.W   R13
						   50447 => x"6D",
						   50448 => x"09",		-- 00c510: 0969             RLC.W   R9
						   50449 => x"69",
						   50450 => x"09",		-- 00c512: 098E             SUB.W   R14,R9
						   50451 => x"8E",
						   50452 => x"04",		-- 00c514: 0428             JLO     (undo_sub)
						   50453 => x"28",
						   50454 => x"1C",		-- 00c516: 1CD3             BIS.W   #1,R12
						   50455 => x"D3",
						   50456 => x"0B",		-- 00c518: 0B5B             RLA.W   R11
						   50457 => x"5B",
						   50458 => x"F8",		-- 00c51a: F82B             JLO     (div_loop_lo)
						   50459 => x"2B",
						   50460 => x"03",		-- 00c51c: 033C             JMP     (process_hi)
						   50461 => x"3C",
						   -- Begin: undo_sub
						   50462 => x"09",		-- 00c51e: 095E             ADD.W   R14,R9
						   50463 => x"5E",
						   50464 => x"0B",		-- 00c520: 0B5B             RLA.W   R11
						   50465 => x"5B",
						   50466 => x"F4",		-- 00c522: F42B             JLO     (div_loop_lo)
						   50467 => x"2B",
						   -- Begin: process_hi
						   50468 => x"1B",		-- 00c524: 1B43             MOV.W   #1,R11
						   50469 => x"43",
						   -- Begin: div_loop_hi
						   50470 => x"0C",		-- 00c526: 0C5C             RLA.W   R12
						   50471 => x"5C",
						   50472 => x"0D",		-- 00c528: 0D6D             RLC.W   R13
						   50473 => x"6D",
						   50474 => x"09",		-- 00c52a: 0969             RLC.W   R9
						   50475 => x"69",
						   50476 => x"0A",		-- 00c52c: 0A6A             RLC.W   R10
						   50477 => x"6A",
						   50478 => x"09",		-- 00c52e: 098E             SUB.W   R14,R9
						   50479 => x"8E",
						   50480 => x"0A",		-- 00c530: 0A7F             SUBC.W  R15,R10
						   50481 => x"7F",
						   50482 => x"04",		-- 00c532: 0428             JLO     (undo_sub_hi)
						   50483 => x"28",
						   50484 => x"1C",		-- 00c534: 1CD3             BIS.W   #1,R12
						   50485 => x"D3",
						   50486 => x"0B",		-- 00c536: 0B5B             RLA.W   R11
						   50487 => x"5B",
						   50488 => x"F6",		-- 00c538: F62B             JLO     (div_loop_hi)
						   50489 => x"2B",
						   50490 => x"04",		-- 00c53a: 043C             JMP     (div_end)
						   50491 => x"3C",
						   -- Begin: undo_sub_hi
						   50492 => x"09",		-- 00c53c: 095E             ADD.W   R14,R9
						   50493 => x"5E",
						   50494 => x"0A",		-- 00c53e: 0A6F             ADDC.W  R15,R10
						   50495 => x"6F",
						   50496 => x"0B",		-- 00c540: 0B5B             RLA.W   R11
						   50497 => x"5B",
						   50498 => x"F1",		-- 00c542: F12B             JLO     (div_loop_hi)
						   50499 => x"2B",
						   -- Begin: div_end
						   50500 => x"0E",		-- 00c544: 0E49             MOV.W   R9,R14
						   50501 => x"49",
						   50502 => x"0F",		-- 00c546: 0F4A             MOV.W   R10,R15
						   50503 => x"4A",
						   50504 => x"39",		-- 00c548: 3941             POP.W   R9
						   50505 => x"41",
						   50506 => x"3A",		-- 00c54a: 3A41             POP.W   R10
						   50507 => x"41",
						   50508 => x"30",		-- 00c54c: 3041             RET     
						   50509 => x"41",
						   -- Begin: atoi
						   50510 => x"0A",		-- 00c54e: 0A12             PUSH    R10
						   50511 => x"12",
						   50512 => x"0B",		-- 00c550: 0B4C             MOV.W   R12,R11
						   50513 => x"4C",
						   50514 => x"0C",		-- 00c552: 0C43             CLR.W   R12
						   50515 => x"43",
						   50516 => x"0B",		-- 00c554: 0B3C             JMP     ($C$L3)
						   50517 => x"3C",
						   50518 => x"3D",		-- 00c556: 3D40             MOV.W   #0x000a,R13
						   50519 => x"40",
						   50520 => x"0A",		-- 00c558: 0A00            
						   50521 => x"00",
						   50522 => x"B0",		-- 00c55a: B012             CALL    #__mspabi_mpyi
						   50523 => x"12",
						   50524 => x"2C",		-- 00c55c: 2CCD            
						   50525 => x"CD",
						   50526 => x"0C",		-- 00c55e: 0C5F             ADD.W   R15,R12
						   50527 => x"5F",
						   50528 => x"3C",		-- 00c560: 3C80             SUB.W   #0x0030,R12
						   50529 => x"80",
						   50530 => x"30",		-- 00c562: 3000            
						   50531 => x"00",
						   50532 => x"1B",		-- 00c564: 1B53             INC.W   R11
						   50533 => x"53",
						   50534 => x"6F",		-- 00c566: 6F4B             MOV.B   @R11,R15
						   50535 => x"4B",
						   50536 => x"12",		-- 00c568: 123C             JMP     ($C$L6)
						   50537 => x"3C",
						   50538 => x"1B",		-- 00c56a: 1B53             INC.W   R11
						   50539 => x"53",
						   50540 => x"6F",		-- 00c56c: 6F4B             MOV.B   @R11,R15
						   50541 => x"4B",
						   50542 => x"4E",		-- 00c56e: 4E4F             MOV.B   R15,R14
						   50543 => x"4F",
						   50544 => x"FE",		-- 00c570: FEB2             BIT.B   #8,0x8515(R14)
						   50545 => x"B2",
						   50546 => x"15",		-- 00c572: 1585            
						   50547 => x"85",
						   50548 => x"FA",		-- 00c574: FA23             JNE     ($C$L2)
						   50549 => x"23",
						   50550 => x"4F",		-- 00c576: 4F4F             MOV.B   R15,R15
						   50551 => x"4F",
						   50552 => x"3F",		-- 00c578: 3F90             CMP.W   #0x002d,R15
						   50553 => x"90",
						   50554 => x"2D",		-- 00c57a: 2D00            
						   50555 => x"00",
						   50556 => x"05",		-- 00c57c: 0524             JEQ     ($C$L4)
						   50557 => x"24",
						   50558 => x"0A",		-- 00c57e: 0A43             CLR.W   R10
						   50559 => x"43",
						   50560 => x"3F",		-- 00c580: 3F90             CMP.W   #0x002b,R15
						   50561 => x"90",
						   50562 => x"2B",		-- 00c582: 2B00            
						   50563 => x"00",
						   50564 => x"04",		-- 00c584: 0420             JNE     ($C$L6)
						   50565 => x"20",
						   50566 => x"01",		-- 00c586: 013C             JMP     ($C$L5)
						   50567 => x"3C",
						   50568 => x"1A",		-- 00c588: 1A43             MOV.W   #1,R10
						   50569 => x"43",
						   50570 => x"1B",		-- 00c58a: 1B53             INC.W   R11
						   50571 => x"53",
						   50572 => x"6F",		-- 00c58c: 6F4B             MOV.B   @R11,R15
						   50573 => x"4B",
						   50574 => x"EF",		-- 00c58e: EFB2             BIT.B   #4,0x8515(R15)
						   50575 => x"B2",
						   50576 => x"15",		-- 00c590: 1585            
						   50577 => x"85",
						   50578 => x"E1",		-- 00c592: E123             JNE     ($C$L1)
						   50579 => x"23",
						   50580 => x"0A",		-- 00c594: 0A93             TST.W   R10
						   50581 => x"93",
						   50582 => x"02",		-- 00c596: 0224             JEQ     ($C$L7)
						   50583 => x"24",
						   50584 => x"3C",		-- 00c598: 3CE3             INV.W   R12
						   50585 => x"E3",
						   50586 => x"1C",		-- 00c59a: 1C53             INC.W   R12
						   50587 => x"53",
						   50588 => x"3A",		-- 00c59c: 3A41             POP.W   R10
						   50589 => x"41",
						   50590 => x"30",		-- 00c59e: 3041             RET     
						   50591 => x"41",
						   -- Begin: _fcpy
						   50592 => x"0A",		-- 00c5a0: 0A12             PUSH    R10
						   50593 => x"12",
						   50594 => x"09",		-- 00c5a2: 0912             PUSH    R9
						   50595 => x"12",
						   50596 => x"08",		-- 00c5a4: 0812             PUSH    R8
						   50597 => x"12",
						   50598 => x"07",		-- 00c5a6: 0712             PUSH    R7
						   50599 => x"12",
						   50600 => x"08",		-- 00c5a8: 084F             MOV.W   R15,R8
						   50601 => x"4F",
						   50602 => x"09",		-- 00c5aa: 094E             MOV.W   R14,R9
						   50603 => x"4E",
						   50604 => x"07",		-- 00c5ac: 074C             MOV.W   R12,R7
						   50605 => x"4C",
						   50606 => x"0D",		-- 00c5ae: 0D59             ADD.W   R9,R13
						   50607 => x"59",
						   50608 => x"1D",		-- 00c5b0: 1D83             DEC.W   R13
						   50609 => x"83",
						   50610 => x"0A",		-- 00c5b2: 0A4D             MOV.W   R13,R10
						   50611 => x"4D",
						   50612 => x"B0",		-- 00c5b4: B012             CALL    #strlen
						   50613 => x"12",
						   50614 => x"BC",		-- 00c5b6: BCCD            
						   50615 => x"CD",
						   50616 => x"19",		-- 00c5b8: 1983             DEC.W   R9
						   50617 => x"83",
						   50618 => x"09",		-- 00c5ba: 0993             TST.W   R9
						   50619 => x"93",
						   50620 => x"16",		-- 00c5bc: 1638             JL      ($C$L149)
						   50621 => x"38",
						   50622 => x"1E",		-- 00c5be: 1E43             MOV.W   #1,R14
						   50623 => x"43",
						   50624 => x"0E",		-- 00c5c0: 0E59             ADD.W   R9,R14
						   50625 => x"59",
						   50626 => x"0A",		-- 00c5c2: 0A93             TST.W   R10
						   50627 => x"93",
						   50628 => x"06",		-- 00c5c4: 0638             JL      ($C$L147)
						   50629 => x"38",
						   50630 => x"0A",		-- 00c5c6: 0A9C             CMP.W   R12,R10
						   50631 => x"9C",
						   50632 => x"04",		-- 00c5c8: 0434             JGE     ($C$L147)
						   50633 => x"34",
						   50634 => x"0F",		-- 00c5ca: 0F4A             MOV.W   R10,R15
						   50635 => x"4A",
						   50636 => x"0F",		-- 00c5cc: 0F57             ADD.W   R7,R15
						   50637 => x"57",
						   50638 => x"6D",		-- 00c5ce: 6D4F             MOV.B   @R15,R13
						   50639 => x"4F",
						   50640 => x"02",		-- 00c5d0: 023C             JMP     ($C$L148)
						   50641 => x"3C",
						   50642 => x"3D",		-- 00c5d2: 3D40             MOV.W   #0x0030,R13
						   50643 => x"40",
						   50644 => x"30",		-- 00c5d4: 3000            
						   50645 => x"00",
						   50646 => x"2B",		-- 00c5d6: 2B48             MOV.W   @R8,R11
						   50647 => x"48",
						   50648 => x"0F",		-- 00c5d8: 0F4B             MOV.W   R11,R15
						   50649 => x"4B",
						   50650 => x"1F",		-- 00c5da: 1F83             DEC.W   R15
						   50651 => x"83",
						   50652 => x"88",		-- 00c5dc: 884F             MOV.W   R15,0x0000(R8)
						   50653 => x"4F",
						   50654 => x"00",		-- 00c5de: 0000            
						   50655 => x"00",
						   50656 => x"CB",		-- 00c5e0: CB4D             MOV.B   R13,0x0000(R11)
						   50657 => x"4D",
						   50658 => x"00",		-- 00c5e2: 0000            
						   50659 => x"00",
						   50660 => x"1A",		-- 00c5e4: 1A83             DEC.W   R10
						   50661 => x"83",
						   50662 => x"1E",		-- 00c5e6: 1E83             DEC.W   R14
						   50663 => x"83",
						   50664 => x"EC",		-- 00c5e8: EC23             JNE     ($C$L146)
						   50665 => x"23",
						   50666 => x"30",		-- 00c5ea: 3040             BR      #__mspabi_func_epilog_4
						   50667 => x"40",
						   50668 => x"A2",		-- 00c5ec: A2CD            
						   50669 => x"CD",
						   -- Begin: __mspabi_srli
						   50670 => x"3D",		-- 00c5ee: 3DF0             AND.W   #0x000f,R13
						   50671 => x"F0",
						   50672 => x"0F",		-- 00c5f0: 0F00            
						   50673 => x"00",
						   50674 => x"3D",		-- 00c5f2: 3DE0             XOR.W   #0x000f,R13
						   50675 => x"E0",
						   50676 => x"0F",		-- 00c5f4: 0F00            
						   50677 => x"00",
						   50678 => x"0D",		-- 00c5f6: 0D5D             RLA.W   R13
						   50679 => x"5D",
						   50680 => x"0D",		-- 00c5f8: 0D5D             RLA.W   R13
						   50681 => x"5D",
						   50682 => x"00",		-- 00c5fa: 005D             ADD.W   R13,PC
						   50683 => x"5D",
						   -- Begin: __mspabi_srli_15
						   50684 => x"12",		-- 00c5fc: 12C3             CLRC    
						   50685 => x"C3",
						   50686 => x"0C",		-- 00c5fe: 0C10             RRC     R12
						   50687 => x"10",
						   -- Begin: __mspabi_srli_14
						   50688 => x"12",		-- 00c600: 12C3             CLRC    
						   50689 => x"C3",
						   50690 => x"0C",		-- 00c602: 0C10             RRC     R12
						   50691 => x"10",
						   -- Begin: __mspabi_srli_13
						   50692 => x"12",		-- 00c604: 12C3             CLRC    
						   50693 => x"C3",
						   50694 => x"0C",		-- 00c606: 0C10             RRC     R12
						   50695 => x"10",
						   -- Begin: __mspabi_srli_12
						   50696 => x"12",		-- 00c608: 12C3             CLRC    
						   50697 => x"C3",
						   50698 => x"0C",		-- 00c60a: 0C10             RRC     R12
						   50699 => x"10",
						   -- Begin: __mspabi_srli_11
						   50700 => x"12",		-- 00c60c: 12C3             CLRC    
						   50701 => x"C3",
						   50702 => x"0C",		-- 00c60e: 0C10             RRC     R12
						   50703 => x"10",
						   -- Begin: __mspabi_srli_10
						   50704 => x"12",		-- 00c610: 12C3             CLRC    
						   50705 => x"C3",
						   50706 => x"0C",		-- 00c612: 0C10             RRC     R12
						   50707 => x"10",
						   -- Begin: __mspabi_srli_9
						   50708 => x"12",		-- 00c614: 12C3             CLRC    
						   50709 => x"C3",
						   50710 => x"0C",		-- 00c616: 0C10             RRC     R12
						   50711 => x"10",
						   -- Begin: __mspabi_srli_8
						   50712 => x"12",		-- 00c618: 12C3             CLRC    
						   50713 => x"C3",
						   50714 => x"0C",		-- 00c61a: 0C10             RRC     R12
						   50715 => x"10",
						   -- Begin: __mspabi_srli_7
						   50716 => x"12",		-- 00c61c: 12C3             CLRC    
						   50717 => x"C3",
						   50718 => x"0C",		-- 00c61e: 0C10             RRC     R12
						   50719 => x"10",
						   -- Begin: __mspabi_srli_6
						   50720 => x"12",		-- 00c620: 12C3             CLRC    
						   50721 => x"C3",
						   50722 => x"0C",		-- 00c622: 0C10             RRC     R12
						   50723 => x"10",
						   -- Begin: __mspabi_srli_5
						   50724 => x"12",		-- 00c624: 12C3             CLRC    
						   50725 => x"C3",
						   50726 => x"0C",		-- 00c626: 0C10             RRC     R12
						   50727 => x"10",
						   -- Begin: __mspabi_srli_4
						   50728 => x"12",		-- 00c628: 12C3             CLRC    
						   50729 => x"C3",
						   50730 => x"0C",		-- 00c62a: 0C10             RRC     R12
						   50731 => x"10",
						   -- Begin: __mspabi_srli_3
						   50732 => x"12",		-- 00c62c: 12C3             CLRC    
						   50733 => x"C3",
						   50734 => x"0C",		-- 00c62e: 0C10             RRC     R12
						   50735 => x"10",
						   -- Begin: __mspabi_srli_2
						   50736 => x"12",		-- 00c630: 12C3             CLRC    
						   50737 => x"C3",
						   50738 => x"0C",		-- 00c632: 0C10             RRC     R12
						   50739 => x"10",
						   -- Begin: __mspabi_srli_1
						   50740 => x"12",		-- 00c634: 12C3             CLRC    
						   50741 => x"C3",
						   50742 => x"0C",		-- 00c636: 0C10             RRC     R12
						   50743 => x"10",
						   50744 => x"30",		-- 00c638: 3041             RET     
						   50745 => x"41",
						   -- Begin: __mspabi_srall
						   50746 => x"07",		-- 00c63a: 0712             PUSH    R7
						   50747 => x"12",
						   50748 => x"07",		-- 00c63c: 074C             MOV.W   R12,R7
						   50749 => x"4C",
						   50750 => x"0D",		-- 00c63e: 0D49             MOV.W   R9,R13
						   50751 => x"49",
						   50752 => x"0E",		-- 00c640: 0E4A             MOV.W   R10,R14
						   50753 => x"4A",
						   50754 => x"0F",		-- 00c642: 0F4B             MOV.W   R11,R15
						   50755 => x"4B",
						   50756 => x"37",		-- 00c644: 3790             CMP.W   #0x0011,R7
						   50757 => x"90",
						   50758 => x"11",		-- 00c646: 1100            
						   50759 => x"00",
						   50760 => x"11",		-- 00c648: 1138             JL      ($C$L2)
						   50761 => x"38",
						   50762 => x"0B",		-- 00c64a: 0B47             MOV.W   R7,R11
						   50763 => x"47",
						   50764 => x"1B",		-- 00c64c: 1B83             DEC.W   R11
						   50765 => x"83",
						   50766 => x"0C",		-- 00c64e: 0C4B             MOV.W   R11,R12
						   50767 => x"4B",
						   50768 => x"B0",		-- 00c650: B012             CALL    #__mspabi_srai_4
						   50769 => x"12",
						   50770 => x"9A",		-- 00c652: 9ACA            
						   50771 => x"CA",
						   50772 => x"3B",		-- 00c654: 3BF0             AND.W   #0xfff0,R11
						   50773 => x"F0",
						   50774 => x"F0",		-- 00c656: F0FF            
						   50775 => x"FF",
						   50776 => x"07",		-- 00c658: 078B             SUB.W   R11,R7
						   50777 => x"8B",
						   50778 => x"08",		-- 00c65a: 084D             MOV.W   R13,R8
						   50779 => x"4D",
						   50780 => x"0D",		-- 00c65c: 0D4E             MOV.W   R14,R13
						   50781 => x"4E",
						   50782 => x"0E",		-- 00c65e: 0E4F             MOV.W   R15,R14
						   50783 => x"4F",
						   50784 => x"3F",		-- 00c660: 3FB0             BIT.W   #0x8000,R15
						   50785 => x"B0",
						   50786 => x"00",		-- 00c662: 0080            
						   50787 => x"80",
						   50788 => x"0F",		-- 00c664: 0F7F             SUBC.W  R15,R15
						   50789 => x"7F",
						   50790 => x"3F",		-- 00c666: 3FE3             INV.W   R15
						   50791 => x"E3",
						   50792 => x"1C",		-- 00c668: 1C83             DEC.W   R12
						   50793 => x"83",
						   50794 => x"F7",		-- 00c66a: F723             JNE     ($C$L1)
						   50795 => x"23",
						   50796 => x"17",		-- 00c66c: 1793             CMP.W   #1,R7
						   50797 => x"93",
						   50798 => x"07",		-- 00c66e: 0738             JL      ($C$L4)
						   50799 => x"38",
						   50800 => x"0C",		-- 00c670: 0C47             MOV.W   R7,R12
						   50801 => x"47",
						   50802 => x"0F",		-- 00c672: 0F11             RRA     R15
						   50803 => x"11",
						   50804 => x"0E",		-- 00c674: 0E10             RRC     R14
						   50805 => x"10",
						   50806 => x"0D",		-- 00c676: 0D10             RRC     R13
						   50807 => x"10",
						   50808 => x"08",		-- 00c678: 0810             RRC     R8
						   50809 => x"10",
						   50810 => x"1C",		-- 00c67a: 1C83             DEC.W   R12
						   50811 => x"83",
						   50812 => x"FA",		-- 00c67c: FA23             JNE     ($C$L3)
						   50813 => x"23",
						   50814 => x"0C",		-- 00c67e: 0C48             MOV.W   R8,R12
						   50815 => x"48",
						   50816 => x"37",		-- 00c680: 3741             POP.W   R7
						   50817 => x"41",
						   50818 => x"30",		-- 00c682: 3041             RET     
						   50819 => x"41",
						   -- Begin: close
						   50820 => x"0A",		-- 00c684: 0A12             PUSH    R10
						   50821 => x"12",
						   50822 => x"0A",		-- 00c686: 0A4C             MOV.W   R12,R10
						   50823 => x"4C",
						   50824 => x"0A",		-- 00c688: 0A93             TST.W   R10
						   50825 => x"93",
						   50826 => x"03",		-- 00c68a: 0338             JL      ($C$L1)
						   50827 => x"38",
						   50828 => x"3A",		-- 00c68c: 3A90             CMP.W   #0x000a,R10
						   50829 => x"90",
						   50830 => x"0A",		-- 00c68e: 0A00            
						   50831 => x"00",
						   50832 => x"02",		-- 00c690: 0238             JL      ($C$L2)
						   50833 => x"38",
						   50834 => x"3A",		-- 00c692: 3A43             MOV.W   #-1,R10
						   50835 => x"43",
						   50836 => x"19",		-- 00c694: 193C             JMP     ($C$L6)
						   50837 => x"3C",
						   50838 => x"92",		-- 00c696: 9212             CALL    &_lock
						   50839 => x"12",
						   50840 => x"F2",		-- 00c698: F220            
						   50841 => x"20",
						   50842 => x"0A",		-- 00c69a: 0A5A             RLA.W   R10
						   50843 => x"5A",
						   50844 => x"0A",		-- 00c69c: 0A5A             RLA.W   R10
						   50845 => x"5A",
						   50846 => x"3A",		-- 00c69e: 3A50             ADD.W   #0x20c6,R10
						   50847 => x"50",
						   50848 => x"C6",		-- 00c6a0: C620            
						   50849 => x"20",
						   50850 => x"2F",		-- 00c6a2: 2F4A             MOV.W   @R10,R15
						   50851 => x"4A",
						   50852 => x"0F",		-- 00c6a4: 0F93             TST.W   R15
						   50853 => x"93",
						   50854 => x"02",		-- 00c6a6: 0220             JNE     ($C$L3)
						   50855 => x"20",
						   50856 => x"3A",		-- 00c6a8: 3A43             MOV.W   #-1,R10
						   50857 => x"43",
						   50858 => x"0C",		-- 00c6aa: 0C3C             JMP     ($C$L5)
						   50859 => x"3C",
						   50860 => x"1C",		-- 00c6ac: 1C4A             MOV.W   0x0002(R10),R12
						   50861 => x"4A",
						   50862 => x"02",		-- 00c6ae: 0200            
						   50863 => x"00",
						   50864 => x"9F",		-- 00c6b0: 9F12             CALL    0x000e(R15)
						   50865 => x"12",
						   50866 => x"0E",		-- 00c6b2: 0E00            
						   50867 => x"00",
						   50868 => x"3C",		-- 00c6b4: 3C93             CMP.W   #-1,R12
						   50869 => x"93",
						   50870 => x"05",		-- 00c6b6: 0524             JEQ     ($C$L4)
						   50871 => x"24",
						   50872 => x"2F",		-- 00c6b8: 2F4A             MOV.W   @R10,R15
						   50873 => x"4A",
						   50874 => x"9F",		-- 00c6ba: 9FC3             BIC.W   #1,0x000a(R15)
						   50875 => x"C3",
						   50876 => x"0A",		-- 00c6bc: 0A00            
						   50877 => x"00",
						   50878 => x"8A",		-- 00c6be: 8A43             CLR.W   0x0000(R10)
						   50879 => x"43",
						   50880 => x"00",		-- 00c6c0: 0000            
						   50881 => x"00",
						   50882 => x"0A",		-- 00c6c2: 0A4C             MOV.W   R12,R10
						   50883 => x"4C",
						   50884 => x"92",		-- 00c6c4: 9212             CALL    &_unlock
						   50885 => x"12",
						   50886 => x"F4",		-- 00c6c6: F420            
						   50887 => x"20",
						   50888 => x"0C",		-- 00c6c8: 0C4A             MOV.W   R10,R12
						   50889 => x"4A",
						   50890 => x"3A",		-- 00c6ca: 3A41             POP.W   R10
						   50891 => x"41",
						   50892 => x"30",		-- 00c6cc: 3041             RET     
						   50893 => x"41",
						   -- Begin: __mspabi_srlll
						   50894 => x"07",		-- 00c6ce: 0712             PUSH    R7
						   50895 => x"12",
						   50896 => x"07",		-- 00c6d0: 074C             MOV.W   R12,R7
						   50897 => x"4C",
						   50898 => x"0D",		-- 00c6d2: 0D49             MOV.W   R9,R13
						   50899 => x"49",
						   50900 => x"0E",		-- 00c6d4: 0E4A             MOV.W   R10,R14
						   50901 => x"4A",
						   50902 => x"0F",		-- 00c6d6: 0F4B             MOV.W   R11,R15
						   50903 => x"4B",
						   50904 => x"37",		-- 00c6d8: 3790             CMP.W   #0x0011,R7
						   50905 => x"90",
						   50906 => x"11",		-- 00c6da: 1100            
						   50907 => x"00",
						   50908 => x"0E",		-- 00c6dc: 0E38             JL      ($C$L2)
						   50909 => x"38",
						   50910 => x"0B",		-- 00c6de: 0B47             MOV.W   R7,R11
						   50911 => x"47",
						   50912 => x"1B",		-- 00c6e0: 1B83             DEC.W   R11
						   50913 => x"83",
						   50914 => x"0C",		-- 00c6e2: 0C4B             MOV.W   R11,R12
						   50915 => x"4B",
						   50916 => x"B0",		-- 00c6e4: B012             CALL    #__mspabi_srai_4
						   50917 => x"12",
						   50918 => x"9A",		-- 00c6e6: 9ACA            
						   50919 => x"CA",
						   50920 => x"3B",		-- 00c6e8: 3BF0             AND.W   #0xfff0,R11
						   50921 => x"F0",
						   50922 => x"F0",		-- 00c6ea: F0FF            
						   50923 => x"FF",
						   50924 => x"07",		-- 00c6ec: 078B             SUB.W   R11,R7
						   50925 => x"8B",
						   50926 => x"08",		-- 00c6ee: 084D             MOV.W   R13,R8
						   50927 => x"4D",
						   50928 => x"0D",		-- 00c6f0: 0D4E             MOV.W   R14,R13
						   50929 => x"4E",
						   50930 => x"0E",		-- 00c6f2: 0E4F             MOV.W   R15,R14
						   50931 => x"4F",
						   50932 => x"0F",		-- 00c6f4: 0F43             CLR.W   R15
						   50933 => x"43",
						   50934 => x"1C",		-- 00c6f6: 1C83             DEC.W   R12
						   50935 => x"83",
						   50936 => x"FA",		-- 00c6f8: FA23             JNE     ($C$L1)
						   50937 => x"23",
						   50938 => x"17",		-- 00c6fa: 1793             CMP.W   #1,R7
						   50939 => x"93",
						   50940 => x"08",		-- 00c6fc: 0838             JL      ($C$L4)
						   50941 => x"38",
						   50942 => x"0C",		-- 00c6fe: 0C47             MOV.W   R7,R12
						   50943 => x"47",
						   50944 => x"12",		-- 00c700: 12C3             CLRC    
						   50945 => x"C3",
						   50946 => x"0F",		-- 00c702: 0F10             RRC     R15
						   50947 => x"10",
						   50948 => x"0E",		-- 00c704: 0E10             RRC     R14
						   50949 => x"10",
						   50950 => x"0D",		-- 00c706: 0D10             RRC     R13
						   50951 => x"10",
						   50952 => x"08",		-- 00c708: 0810             RRC     R8
						   50953 => x"10",
						   50954 => x"1C",		-- 00c70a: 1C83             DEC.W   R12
						   50955 => x"83",
						   50956 => x"F9",		-- 00c70c: F923             JNE     ($C$L3)
						   50957 => x"23",
						   50958 => x"0C",		-- 00c70e: 0C48             MOV.W   R8,R12
						   50959 => x"48",
						   50960 => x"37",		-- 00c710: 3741             POP.W   R7
						   50961 => x"41",
						   50962 => x"30",		-- 00c712: 3041             RET     
						   50963 => x"41",
						   -- Begin: HOSTclose
						   50964 => x"0A",		-- 00c714: 0A12             PUSH    R10
						   50965 => x"12",
						   50966 => x"0A",		-- 00c716: 0A4C             MOV.W   R12,R10
						   50967 => x"4C",
						   50968 => x"92",		-- 00c718: 9212             CALL    &_lock
						   50969 => x"12",
						   50970 => x"F2",		-- 00c71a: F220            
						   50971 => x"20",
						   50972 => x"C2",		-- 00c71c: C24A             MOV.B   R10,&parmbuf
						   50973 => x"4A",
						   50974 => x"9E",		-- 00c71e: 9E21            
						   50975 => x"21",
						   50976 => x"8A",		-- 00c720: 8A10             SWPB    R10
						   50977 => x"10",
						   50978 => x"8A",		-- 00c722: 8A11             SXT     R10
						   50979 => x"11",
						   50980 => x"C2",		-- 00c724: C24A             MOV.B   R10,&0x219f
						   50981 => x"4A",
						   50982 => x"9F",		-- 00c726: 9F21            
						   50983 => x"21",
						   50984 => x"7C",		-- 00c728: 7C40             MOV.B   #0x00f1,R12
						   50985 => x"40",
						   50986 => x"F1",		-- 00c72a: F100            
						   50987 => x"00",
						   50988 => x"3D",		-- 00c72c: 3D40             MOV.W   #0x219e,R13
						   50989 => x"40",
						   50990 => x"9E",		-- 00c72e: 9E21            
						   50991 => x"21",
						   50992 => x"0E",		-- 00c730: 0E43             CLR.W   R14
						   50993 => x"43",
						   50994 => x"0F",		-- 00c732: 0F43             CLR.W   R15
						   50995 => x"43",
						   50996 => x"B0",		-- 00c734: B012             CALL    #__TI_writemsg
						   50997 => x"12",
						   50998 => x"C2",		-- 00c736: C2C9            
						   50999 => x"C9",
						   51000 => x"3C",		-- 00c738: 3C40             MOV.W   #0x219e,R12
						   51001 => x"40",
						   51002 => x"9E",		-- 00c73a: 9E21            
						   51003 => x"21",
						   51004 => x"0D",		-- 00c73c: 0D43             CLR.W   R13
						   51005 => x"43",
						   51006 => x"B0",		-- 00c73e: B012             CALL    #__TI_readmsg
						   51007 => x"12",
						   51008 => x"4C",		-- 00c740: 4CCA            
						   51009 => x"CA",
						   51010 => x"5F",		-- 00c742: 5F42             MOV.B   &parmbuf,R15
						   51011 => x"42",
						   51012 => x"9E",		-- 00c744: 9E21            
						   51013 => x"21",
						   51014 => x"5A",		-- 00c746: 5A42             MOV.B   &0x219f,R10
						   51015 => x"42",
						   51016 => x"9F",		-- 00c748: 9F21            
						   51017 => x"21",
						   51018 => x"8A",		-- 00c74a: 8A10             SWPB    R10
						   51019 => x"10",
						   51020 => x"0A",		-- 00c74c: 0A5F             ADD.W   R15,R10
						   51021 => x"5F",
						   51022 => x"92",		-- 00c74e: 9212             CALL    &_unlock
						   51023 => x"12",
						   51024 => x"F4",		-- 00c750: F420            
						   51025 => x"20",
						   51026 => x"0C",		-- 00c752: 0C4A             MOV.W   R10,R12
						   51027 => x"4A",
						   51028 => x"3A",		-- 00c754: 3A41             POP.W   R10
						   51029 => x"41",
						   51030 => x"30",		-- 00c756: 3041             RET     
						   51031 => x"41",
						   -- Begin: __mspabi_sllll
						   51032 => x"07",		-- 00c758: 0712             PUSH    R7
						   51033 => x"12",
						   51034 => x"07",		-- 00c75a: 074C             MOV.W   R12,R7
						   51035 => x"4C",
						   51036 => x"0D",		-- 00c75c: 0D49             MOV.W   R9,R13
						   51037 => x"49",
						   51038 => x"0E",		-- 00c75e: 0E4A             MOV.W   R10,R14
						   51039 => x"4A",
						   51040 => x"0F",		-- 00c760: 0F4B             MOV.W   R11,R15
						   51041 => x"4B",
						   51042 => x"37",		-- 00c762: 3790             CMP.W   #0x0011,R7
						   51043 => x"90",
						   51044 => x"11",		-- 00c764: 1100            
						   51045 => x"00",
						   51046 => x"0E",		-- 00c766: 0E38             JL      ($C$L2)
						   51047 => x"38",
						   51048 => x"0F",		-- 00c768: 0F47             MOV.W   R7,R15
						   51049 => x"47",
						   51050 => x"1F",		-- 00c76a: 1F83             DEC.W   R15
						   51051 => x"83",
						   51052 => x"0C",		-- 00c76c: 0C4F             MOV.W   R15,R12
						   51053 => x"4F",
						   51054 => x"B0",		-- 00c76e: B012             CALL    #__mspabi_srai_4
						   51055 => x"12",
						   51056 => x"9A",		-- 00c770: 9ACA            
						   51057 => x"CA",
						   51058 => x"3F",		-- 00c772: 3FF0             AND.W   #0xfff0,R15
						   51059 => x"F0",
						   51060 => x"F0",		-- 00c774: F0FF            
						   51061 => x"FF",
						   51062 => x"07",		-- 00c776: 078F             SUB.W   R15,R7
						   51063 => x"8F",
						   51064 => x"0F",		-- 00c778: 0F4E             MOV.W   R14,R15
						   51065 => x"4E",
						   51066 => x"0E",		-- 00c77a: 0E4D             MOV.W   R13,R14
						   51067 => x"4D",
						   51068 => x"0D",		-- 00c77c: 0D48             MOV.W   R8,R13
						   51069 => x"48",
						   51070 => x"08",		-- 00c77e: 0843             CLR.W   R8
						   51071 => x"43",
						   51072 => x"1C",		-- 00c780: 1C83             DEC.W   R12
						   51073 => x"83",
						   51074 => x"FA",		-- 00c782: FA23             JNE     ($C$L1)
						   51075 => x"23",
						   51076 => x"17",		-- 00c784: 1793             CMP.W   #1,R7
						   51077 => x"93",
						   51078 => x"07",		-- 00c786: 0738             JL      ($C$L4)
						   51079 => x"38",
						   51080 => x"0C",		-- 00c788: 0C47             MOV.W   R7,R12
						   51081 => x"47",
						   51082 => x"08",		-- 00c78a: 0858             RLA.W   R8
						   51083 => x"58",
						   51084 => x"0D",		-- 00c78c: 0D6D             RLC.W   R13
						   51085 => x"6D",
						   51086 => x"0E",		-- 00c78e: 0E6E             RLC.W   R14
						   51087 => x"6E",
						   51088 => x"0F",		-- 00c790: 0F6F             RLC.W   R15
						   51089 => x"6F",
						   51090 => x"1C",		-- 00c792: 1C83             DEC.W   R12
						   51091 => x"83",
						   51092 => x"FA",		-- 00c794: FA23             JNE     ($C$L3)
						   51093 => x"23",
						   51094 => x"0C",		-- 00c796: 0C48             MOV.W   R8,R12
						   51095 => x"48",
						   51096 => x"37",		-- 00c798: 3741             POP.W   R7
						   51097 => x"41",
						   51098 => x"30",		-- 00c79a: 3041             RET     
						   51099 => x"41",
						   -- Begin: exit
						   51100 => x"0A",		-- 00c79c: 0A12             PUSH    R10
						   51101 => x"12",
						   51102 => x"0A",		-- 00c79e: 0A4C             MOV.W   R12,R10
						   51103 => x"4C",
						   51104 => x"82",		-- 00c7a0: 8293             TST.W   &__TI_enable_exit_profile_output
						   51105 => x"93",
						   51106 => x"FA",		-- 00c7a2: FA20            
						   51107 => x"20",
						   51108 => x"0A",		-- 00c7a4: 0A24             JEQ     ($C$L3)
						   51109 => x"24",
						   51110 => x"3E",		-- 00c7a6: 3E40             MOV.W   #0xffff,R14
						   51111 => x"40",
						   51112 => x"FF",		-- 00c7a8: FFFF            
						   51113 => x"FF",
						   51114 => x"3F",		-- 00c7aa: 3F40             MOV.W   #0xffff,R15
						   51115 => x"40",
						   51116 => x"FF",		-- 00c7ac: FFFF            
						   51117 => x"FF",
						   51118 => x"3F",		-- 00c7ae: 3F93             CMP.W   #-1,R15
						   51119 => x"93",
						   51120 => x"02",		-- 00c7b0: 0220             JNE     ($C$L2)
						   51121 => x"20",
						   51122 => x"3E",		-- 00c7b2: 3E93             CMP.W   #-1,R14
						   51123 => x"93",
						   51124 => x"02",		-- 00c7b4: 0224             JEQ     ($C$L3)
						   51125 => x"24",
						   51126 => x"B0",		-- 00c7b6: B012             CALL    #0xffff
						   51127 => x"12",
						   51128 => x"FF",		-- 00c7b8: FFFF            
						   51129 => x"FF",
						   51130 => x"92",		-- 00c7ba: 9212             CALL    &_lock
						   51131 => x"12",
						   51132 => x"F2",		-- 00c7bc: F220            
						   51133 => x"20",
						   51134 => x"82",		-- 00c7be: 8293             TST.W   &__TI_dtors_ptr
						   51135 => x"93",
						   51136 => x"F0",		-- 00c7c0: F020            
						   51137 => x"20",
						   51138 => x"03",		-- 00c7c2: 0324             JEQ     ($C$L4)
						   51139 => x"24",
						   51140 => x"0C",		-- 00c7c4: 0C4A             MOV.W   R10,R12
						   51141 => x"4A",
						   51142 => x"92",		-- 00c7c6: 9212             CALL    &__TI_dtors_ptr
						   51143 => x"12",
						   51144 => x"F0",		-- 00c7c8: F020            
						   51145 => x"20",
						   51146 => x"82",		-- 00c7ca: 8293             TST.W   &__TI_cleanup_ptr
						   51147 => x"93",
						   51148 => x"EE",		-- 00c7cc: EE20            
						   51149 => x"20",
						   51150 => x"02",		-- 00c7ce: 0224             JEQ     ($C$L5)
						   51151 => x"24",
						   51152 => x"92",		-- 00c7d0: 9212             CALL    &__TI_cleanup_ptr
						   51153 => x"12",
						   51154 => x"EE",		-- 00c7d2: EE20            
						   51155 => x"20",
						   51156 => x"92",		-- 00c7d4: 9212             CALL    &_unlock
						   51157 => x"12",
						   51158 => x"F4",		-- 00c7d6: F420            
						   51159 => x"20",
						   51160 => x"B0",		-- 00c7d8: B012             CALL    #abort
						   51161 => x"12",
						   51162 => x"FA",		-- 00c7da: FACD            
						   51163 => x"CD",
						   51164 => x"3A",		-- 00c7dc: 3A41             POP.W   R10
						   51165 => x"41",
						   51166 => x"30",		-- 00c7de: 3041             RET     
						   51167 => x"41",
						   -- Begin: __TI_auto_init_nobinit_nopinit
						   51168 => x"0A",		-- 00c7e0: 0A12             PUSH    R10
						   51169 => x"12",
						   51170 => x"09",		-- 00c7e2: 0912             PUSH    R9
						   51171 => x"12",
						   51172 => x"3F",		-- 00c7e4: 3F40             MOV.W   #0x8502,R15
						   51173 => x"40",
						   51174 => x"02",		-- 00c7e6: 0285            
						   51175 => x"85",
						   51176 => x"3F",		-- 00c7e8: 3F90             CMP.W   #0x8508,R15
						   51177 => x"90",
						   51178 => x"08",		-- 00c7ea: 0885            
						   51179 => x"85",
						   51180 => x"16",		-- 00c7ec: 1624             JEQ     ($C$L22)
						   51181 => x"24",
						   51182 => x"3F",		-- 00c7ee: 3F40             MOV.W   #0x850c,R15
						   51183 => x"40",
						   51184 => x"0C",		-- 00c7f0: 0C85            
						   51185 => x"85",
						   51186 => x"3F",		-- 00c7f2: 3F90             CMP.W   #0x8514,R15
						   51187 => x"90",
						   51188 => x"14",		-- 00c7f4: 1485            
						   51189 => x"85",
						   51190 => x"11",		-- 00c7f6: 1124             JEQ     ($C$L22)
						   51191 => x"24",
						   51192 => x"3A",		-- 00c7f8: 3A40             MOV.W   #0x8514,R10
						   51193 => x"40",
						   51194 => x"14",		-- 00c7fa: 1485            
						   51195 => x"85",
						   51196 => x"3A",		-- 00c7fc: 3A80             SUB.W   #0x850c,R10
						   51197 => x"80",
						   51198 => x"0C",		-- 00c7fe: 0C85            
						   51199 => x"85",
						   51200 => x"0A",		-- 00c800: 0A11             RRA     R10
						   51201 => x"11",
						   51202 => x"0A",		-- 00c802: 0A11             RRA     R10
						   51203 => x"11",
						   51204 => x"39",		-- 00c804: 3940             MOV.W   #0x850c,R9
						   51205 => x"40",
						   51206 => x"0C",		-- 00c806: 0C85            
						   51207 => x"85",
						   51208 => x"3C",		-- 00c808: 3C49             MOV.W   @R9+,R12
						   51209 => x"49",
						   51210 => x"7F",		-- 00c80a: 7F4C             MOV.B   @R12+,R15
						   51211 => x"4C",
						   51212 => x"0F",		-- 00c80c: 0F5F             RLA.W   R15
						   51213 => x"5F",
						   51214 => x"1F",		-- 00c80e: 1F4F             MOV.W   0x8502(R15),R15
						   51215 => x"4F",
						   51216 => x"02",		-- 00c810: 0285            
						   51217 => x"85",
						   51218 => x"3D",		-- 00c812: 3D49             MOV.W   @R9+,R13
						   51219 => x"49",
						   51220 => x"8F",		-- 00c814: 8F12             CALL    R15
						   51221 => x"12",
						   51222 => x"1A",		-- 00c816: 1A83             DEC.W   R10
						   51223 => x"83",
						   51224 => x"F7",		-- 00c818: F723             JNE     ($C$L21)
						   51225 => x"23",
						   51226 => x"B0",		-- 00c81a: B012             CALL    #_system_post_cinit
						   51227 => x"12",
						   51228 => x"0A",		-- 00c81c: 0ACE            
						   51229 => x"CE",
						   51230 => x"30",		-- 00c81e: 3040             BR      #__mspabi_func_epilog_2
						   51231 => x"40",
						   51232 => x"A6",		-- 00c820: A6CD            
						   51233 => x"CD",
						   -- Begin: HOSTunlink
						   51234 => x"0A",		-- 00c822: 0A12             PUSH    R10
						   51235 => x"12",
						   51236 => x"0A",		-- 00c824: 0A4C             MOV.W   R12,R10
						   51237 => x"4C",
						   51238 => x"92",		-- 00c826: 9212             CALL    &_lock
						   51239 => x"12",
						   51240 => x"F2",		-- 00c828: F220            
						   51241 => x"20",
						   51242 => x"0C",		-- 00c82a: 0C4A             MOV.W   R10,R12
						   51243 => x"4A",
						   51244 => x"B0",		-- 00c82c: B012             CALL    #strlen
						   51245 => x"12",
						   51246 => x"BC",		-- 00c82e: BCCD            
						   51247 => x"CD",
						   51248 => x"1F",		-- 00c830: 1F43             MOV.W   #1,R15
						   51249 => x"43",
						   51250 => x"0F",		-- 00c832: 0F5C             ADD.W   R12,R15
						   51251 => x"5C",
						   51252 => x"7C",		-- 00c834: 7C40             MOV.B   #0x00f5,R12
						   51253 => x"40",
						   51254 => x"F5",		-- 00c836: F500            
						   51255 => x"00",
						   51256 => x"3D",		-- 00c838: 3D40             MOV.W   #0x219e,R13
						   51257 => x"40",
						   51258 => x"9E",		-- 00c83a: 9E21            
						   51259 => x"21",
						   51260 => x"0E",		-- 00c83c: 0E4A             MOV.W   R10,R14
						   51261 => x"4A",
						   51262 => x"B0",		-- 00c83e: B012             CALL    #__TI_writemsg
						   51263 => x"12",
						   51264 => x"C2",		-- 00c840: C2C9            
						   51265 => x"C9",
						   51266 => x"3C",		-- 00c842: 3C40             MOV.W   #0x219e,R12
						   51267 => x"40",
						   51268 => x"9E",		-- 00c844: 9E21            
						   51269 => x"21",
						   51270 => x"0D",		-- 00c846: 0D43             CLR.W   R13
						   51271 => x"43",
						   51272 => x"B0",		-- 00c848: B012             CALL    #__TI_readmsg
						   51273 => x"12",
						   51274 => x"4C",		-- 00c84a: 4CCA            
						   51275 => x"CA",
						   51276 => x"5F",		-- 00c84c: 5F42             MOV.B   &parmbuf,R15
						   51277 => x"42",
						   51278 => x"9E",		-- 00c84e: 9E21            
						   51279 => x"21",
						   51280 => x"5A",		-- 00c850: 5A42             MOV.B   &0x219f,R10
						   51281 => x"42",
						   51282 => x"9F",		-- 00c852: 9F21            
						   51283 => x"21",
						   51284 => x"8A",		-- 00c854: 8A10             SWPB    R10
						   51285 => x"10",
						   51286 => x"0A",		-- 00c856: 0A5F             ADD.W   R15,R10
						   51287 => x"5F",
						   51288 => x"92",		-- 00c858: 9212             CALL    &_unlock
						   51289 => x"12",
						   51290 => x"F4",		-- 00c85a: F420            
						   51291 => x"20",
						   51292 => x"0C",		-- 00c85c: 0C4A             MOV.W   R10,R12
						   51293 => x"4A",
						   51294 => x"3A",		-- 00c85e: 3A41             POP.W   R10
						   51295 => x"41",
						   51296 => x"30",		-- 00c860: 3041             RET     
						   51297 => x"41",
						   -- Begin: __mspabi_divli
						   -- Begin: __mspabi_remli
						   51298 => x"0A",		-- 00c862: 0A12             PUSH    R10
						   51299 => x"12",
						   51300 => x"0A",		-- 00c864: 0A43             CLR.W   R10
						   51301 => x"43",
						   51302 => x"0F",		-- 00c866: 0F93             TST.W   R15
						   51303 => x"93",
						   51304 => x"05",		-- 00c868: 0534             JGE     (dvd_sign)
						   51305 => x"34",
						   51306 => x"3E",		-- 00c86a: 3EE3             INV.W   R14
						   51307 => x"E3",
						   51308 => x"3F",		-- 00c86c: 3FE3             INV.W   R15
						   51309 => x"E3",
						   51310 => x"1E",		-- 00c86e: 1E53             INC.W   R14
						   51311 => x"53",
						   51312 => x"0F",		-- 00c870: 0F63             ADC.W   R15
						   51313 => x"63",
						   51314 => x"1A",		-- 00c872: 1AD3             BIS.W   #1,R10
						   51315 => x"D3",
						   -- Begin: dvd_sign
						   51316 => x"0D",		-- 00c874: 0D93             TST.W   R13
						   51317 => x"93",
						   51318 => x"05",		-- 00c876: 0534             JGE     (perform_divide)
						   51319 => x"34",
						   51320 => x"3C",		-- 00c878: 3CE3             INV.W   R12
						   51321 => x"E3",
						   51322 => x"3D",		-- 00c87a: 3DE3             INV.W   R13
						   51323 => x"E3",
						   51324 => x"1C",		-- 00c87c: 1C53             INC.W   R12
						   51325 => x"53",
						   51326 => x"0D",		-- 00c87e: 0D63             ADC.W   R13
						   51327 => x"63",
						   51328 => x"3A",		-- 00c880: 3AE3             INV.W   R10
						   51329 => x"E3",
						   -- Begin: perform_divide
						   51330 => x"B0",		-- 00c882: B012             CALL    #__mspabi_divul
						   51331 => x"12",
						   51332 => x"F6",		-- 00c884: F6C4            
						   51333 => x"C4",
						   51334 => x"1A",		-- 00c886: 1AB3             BIT.W   #1,R10
						   51335 => x"B3",
						   51336 => x"04",		-- 00c888: 0424             JEQ     (rem_sign)
						   51337 => x"24",
						   51338 => x"3C",		-- 00c88a: 3CE3             INV.W   R12
						   51339 => x"E3",
						   51340 => x"3D",		-- 00c88c: 3DE3             INV.W   R13
						   51341 => x"E3",
						   51342 => x"1C",		-- 00c88e: 1C53             INC.W   R12
						   51343 => x"53",
						   51344 => x"0D",		-- 00c890: 0D63             ADC.W   R13
						   51345 => x"63",
						   -- Begin: rem_sign
						   51346 => x"2A",		-- 00c892: 2AB3             BIT.W   #2,R10
						   51347 => x"B3",
						   51348 => x"04",		-- 00c894: 0424             JEQ     (div_exit)
						   51349 => x"24",
						   51350 => x"3E",		-- 00c896: 3EE3             INV.W   R14
						   51351 => x"E3",
						   51352 => x"3F",		-- 00c898: 3FE3             INV.W   R15
						   51353 => x"E3",
						   51354 => x"1E",		-- 00c89a: 1E53             INC.W   R14
						   51355 => x"53",
						   51356 => x"0F",		-- 00c89c: 0F63             ADC.W   R15
						   51357 => x"63",
						   -- Begin: div_exit
						   51358 => x"3A",		-- 00c89e: 3A41             POP.W   R10
						   51359 => x"41",
						   51360 => x"30",		-- 00c8a0: 3041             RET     
						   51361 => x"41",
						   -- Begin: __mspabi_sral_15
						   51362 => x"0D",		-- 00c8a2: 0D11             RRA     R13
						   51363 => x"11",
						   51364 => x"0C",		-- 00c8a4: 0C10             RRC     R12
						   51365 => x"10",
						   -- Begin: __mspabi_sral_14
						   51366 => x"0D",		-- 00c8a6: 0D11             RRA     R13
						   51367 => x"11",
						   51368 => x"0C",		-- 00c8a8: 0C10             RRC     R12
						   51369 => x"10",
						   -- Begin: __mspabi_sral_13
						   51370 => x"0D",		-- 00c8aa: 0D11             RRA     R13
						   51371 => x"11",
						   51372 => x"0C",		-- 00c8ac: 0C10             RRC     R12
						   51373 => x"10",
						   -- Begin: __mspabi_sral_12
						   51374 => x"0D",		-- 00c8ae: 0D11             RRA     R13
						   51375 => x"11",
						   51376 => x"0C",		-- 00c8b0: 0C10             RRC     R12
						   51377 => x"10",
						   -- Begin: __mspabi_sral_11
						   51378 => x"0D",		-- 00c8b2: 0D11             RRA     R13
						   51379 => x"11",
						   51380 => x"0C",		-- 00c8b4: 0C10             RRC     R12
						   51381 => x"10",
						   -- Begin: __mspabi_sral_10
						   51382 => x"0D",		-- 00c8b6: 0D11             RRA     R13
						   51383 => x"11",
						   51384 => x"0C",		-- 00c8b8: 0C10             RRC     R12
						   51385 => x"10",
						   -- Begin: __mspabi_sral_9
						   51386 => x"0D",		-- 00c8ba: 0D11             RRA     R13
						   51387 => x"11",
						   51388 => x"0C",		-- 00c8bc: 0C10             RRC     R12
						   51389 => x"10",
						   -- Begin: __mspabi_sral_8
						   51390 => x"0D",		-- 00c8be: 0D11             RRA     R13
						   51391 => x"11",
						   51392 => x"0C",		-- 00c8c0: 0C10             RRC     R12
						   51393 => x"10",
						   -- Begin: __mspabi_sral_7
						   51394 => x"0D",		-- 00c8c2: 0D11             RRA     R13
						   51395 => x"11",
						   51396 => x"0C",		-- 00c8c4: 0C10             RRC     R12
						   51397 => x"10",
						   -- Begin: __mspabi_sral_6
						   51398 => x"0D",		-- 00c8c6: 0D11             RRA     R13
						   51399 => x"11",
						   51400 => x"0C",		-- 00c8c8: 0C10             RRC     R12
						   51401 => x"10",
						   -- Begin: __mspabi_sral_5
						   51402 => x"0D",		-- 00c8ca: 0D11             RRA     R13
						   51403 => x"11",
						   51404 => x"0C",		-- 00c8cc: 0C10             RRC     R12
						   51405 => x"10",
						   -- Begin: __mspabi_sral_4
						   51406 => x"0D",		-- 00c8ce: 0D11             RRA     R13
						   51407 => x"11",
						   51408 => x"0C",		-- 00c8d0: 0C10             RRC     R12
						   51409 => x"10",
						   -- Begin: __mspabi_sral_3
						   51410 => x"0D",		-- 00c8d2: 0D11             RRA     R13
						   51411 => x"11",
						   51412 => x"0C",		-- 00c8d4: 0C10             RRC     R12
						   51413 => x"10",
						   -- Begin: __mspabi_sral_2
						   51414 => x"0D",		-- 00c8d6: 0D11             RRA     R13
						   51415 => x"11",
						   51416 => x"0C",		-- 00c8d8: 0C10             RRC     R12
						   51417 => x"10",
						   -- Begin: __mspabi_sral_1
						   51418 => x"0D",		-- 00c8da: 0D11             RRA     R13
						   51419 => x"11",
						   51420 => x"0C",		-- 00c8dc: 0C10             RRC     R12
						   51421 => x"10",
						   51422 => x"30",		-- 00c8de: 3041             RET     
						   51423 => x"41",
						   -- Begin: __mspabi_slll_15
						   51424 => x"0C",		-- 00c8e0: 0C5C             RLA.W   R12
						   51425 => x"5C",
						   51426 => x"0D",		-- 00c8e2: 0D6D             RLC.W   R13
						   51427 => x"6D",
						   -- Begin: __mspabi_slll_14
						   51428 => x"0C",		-- 00c8e4: 0C5C             RLA.W   R12
						   51429 => x"5C",
						   51430 => x"0D",		-- 00c8e6: 0D6D             RLC.W   R13
						   51431 => x"6D",
						   -- Begin: __mspabi_slll_13
						   51432 => x"0C",		-- 00c8e8: 0C5C             RLA.W   R12
						   51433 => x"5C",
						   51434 => x"0D",		-- 00c8ea: 0D6D             RLC.W   R13
						   51435 => x"6D",
						   -- Begin: __mspabi_slll_12
						   51436 => x"0C",		-- 00c8ec: 0C5C             RLA.W   R12
						   51437 => x"5C",
						   51438 => x"0D",		-- 00c8ee: 0D6D             RLC.W   R13
						   51439 => x"6D",
						   -- Begin: __mspabi_slll_11
						   51440 => x"0C",		-- 00c8f0: 0C5C             RLA.W   R12
						   51441 => x"5C",
						   51442 => x"0D",		-- 00c8f2: 0D6D             RLC.W   R13
						   51443 => x"6D",
						   -- Begin: __mspabi_slll_10
						   51444 => x"0C",		-- 00c8f4: 0C5C             RLA.W   R12
						   51445 => x"5C",
						   51446 => x"0D",		-- 00c8f6: 0D6D             RLC.W   R13
						   51447 => x"6D",
						   -- Begin: __mspabi_slll_9
						   51448 => x"0C",		-- 00c8f8: 0C5C             RLA.W   R12
						   51449 => x"5C",
						   51450 => x"0D",		-- 00c8fa: 0D6D             RLC.W   R13
						   51451 => x"6D",
						   -- Begin: __mspabi_slll_8
						   51452 => x"0C",		-- 00c8fc: 0C5C             RLA.W   R12
						   51453 => x"5C",
						   51454 => x"0D",		-- 00c8fe: 0D6D             RLC.W   R13
						   51455 => x"6D",
						   -- Begin: __mspabi_slll_7
						   51456 => x"0C",		-- 00c900: 0C5C             RLA.W   R12
						   51457 => x"5C",
						   51458 => x"0D",		-- 00c902: 0D6D             RLC.W   R13
						   51459 => x"6D",
						   -- Begin: __mspabi_slll_6
						   51460 => x"0C",		-- 00c904: 0C5C             RLA.W   R12
						   51461 => x"5C",
						   51462 => x"0D",		-- 00c906: 0D6D             RLC.W   R13
						   51463 => x"6D",
						   -- Begin: __mspabi_slll_5
						   51464 => x"0C",		-- 00c908: 0C5C             RLA.W   R12
						   51465 => x"5C",
						   51466 => x"0D",		-- 00c90a: 0D6D             RLC.W   R13
						   51467 => x"6D",
						   -- Begin: __mspabi_slll_4
						   51468 => x"0C",		-- 00c90c: 0C5C             RLA.W   R12
						   51469 => x"5C",
						   51470 => x"0D",		-- 00c90e: 0D6D             RLC.W   R13
						   51471 => x"6D",
						   -- Begin: __mspabi_slll_3
						   51472 => x"0C",		-- 00c910: 0C5C             RLA.W   R12
						   51473 => x"5C",
						   51474 => x"0D",		-- 00c912: 0D6D             RLC.W   R13
						   51475 => x"6D",
						   -- Begin: __mspabi_slll_2
						   51476 => x"0C",		-- 00c914: 0C5C             RLA.W   R12
						   51477 => x"5C",
						   51478 => x"0D",		-- 00c916: 0D6D             RLC.W   R13
						   51479 => x"6D",
						   -- Begin: __mspabi_slll_1
						   51480 => x"0C",		-- 00c918: 0C5C             RLA.W   R12
						   51481 => x"5C",
						   51482 => x"0D",		-- 00c91a: 0D6D             RLC.W   R13
						   51483 => x"6D",
						   51484 => x"30",		-- 00c91c: 3041             RET     
						   51485 => x"41",
						   -- Begin: printf
						   51486 => x"0A",		-- 00c91e: 0A12             PUSH    R10
						   51487 => x"12",
						   51488 => x"21",		-- 00c920: 2183             DECD.W  SP
						   51489 => x"83",
						   51490 => x"92",		-- 00c922: 9212             CALL    &_lock
						   51491 => x"12",
						   51492 => x"F2",		-- 00c924: F220            
						   51493 => x"20",
						   51494 => x"B2",		-- 00c926: B293             CMP.W   #-1,&0x200c
						   51495 => x"93",
						   51496 => x"0C",		-- 00c928: 0C20            
						   51497 => x"20",
						   51498 => x"02",		-- 00c92a: 0220             JNE     ($C$L1)
						   51499 => x"20",
						   51500 => x"3A",		-- 00c92c: 3A43             MOV.W   #-1,R10
						   51501 => x"43",
						   51502 => x"0F",		-- 00c92e: 0F3C             JMP     ($C$L2)
						   51503 => x"3C",
						   51504 => x"B1",		-- 00c930: B140             MOV.W   #0xce00,0x0000(SP)
						   51505 => x"40",
						   51506 => x"00",		-- 00c932: 00CE            
						   51507 => x"CE",
						   51508 => x"00",		-- 00c934: 0000            
						   51509 => x"00",
						   51510 => x"0D",		-- 00c936: 0D41             MOV.W   SP,R13
						   51511 => x"41",
						   51512 => x"3D",		-- 00c938: 3D52             ADD.W   #8,R13
						   51513 => x"52",
						   51514 => x"3E",		-- 00c93a: 3E40             MOV.W   #0x200c,R14
						   51515 => x"40",
						   51516 => x"0C",		-- 00c93c: 0C20            
						   51517 => x"20",
						   51518 => x"0C",		-- 00c93e: 0C41             MOV.W   SP,R12
						   51519 => x"41",
						   51520 => x"3C",		-- 00c940: 3C50             ADD.W   #0x0006,R12
						   51521 => x"50",
						   51522 => x"06",		-- 00c942: 0600            
						   51523 => x"00",
						   51524 => x"3F",		-- 00c944: 3F40             MOV.W   #0xcdf4,R15
						   51525 => x"40",
						   51526 => x"F4",		-- 00c946: F4CD            
						   51527 => x"CD",
						   51528 => x"B0",		-- 00c948: B012             CALL    #__TI_printfi
						   51529 => x"12",
						   51530 => x"32",		-- 00c94a: 3298            
						   51531 => x"98",
						   51532 => x"0A",		-- 00c94c: 0A4C             MOV.W   R12,R10
						   51533 => x"4C",
						   51534 => x"92",		-- 00c94e: 9212             CALL    &_unlock
						   51535 => x"12",
						   51536 => x"F4",		-- 00c950: F420            
						   51537 => x"20",
						   51538 => x"0C",		-- 00c952: 0C4A             MOV.W   R10,R12
						   51539 => x"4A",
						   51540 => x"21",		-- 00c954: 2153             INCD.W  SP
						   51541 => x"53",
						   51542 => x"3A",		-- 00c956: 3A41             POP.W   R10
						   51543 => x"41",
						   51544 => x"30",		-- 00c958: 3041             RET     
						   51545 => x"41",
						   -- Begin: __TI_cleanup
						   51546 => x"0A",		-- 00c95a: 0A12             PUSH    R10
						   51547 => x"12",
						   51548 => x"09",		-- 00c95c: 0912             PUSH    R9
						   51549 => x"12",
						   51550 => x"3C",		-- 00c95e: 3C40             MOV.W   #0x2000,R12
						   51551 => x"40",
						   51552 => x"00",		-- 00c960: 0020            
						   51553 => x"20",
						   51554 => x"B0",		-- 00c962: B012             CALL    #__TI_closefile
						   51555 => x"12",
						   51556 => x"36",		-- 00c964: 36C0            
						   51557 => x"C0",
						   51558 => x"A2",		-- 00c966: A293             CMP.W   #2,&__TI_ft_end
						   51559 => x"93",
						   51560 => x"F6",		-- 00c968: F620            
						   51561 => x"20",
						   51562 => x"0F",		-- 00c96a: 0F38             JL      ($C$L37)
						   51563 => x"38",
						   51564 => x"3A",		-- 00c96c: 3A40             MOV.W   #0x200c,R10
						   51565 => x"40",
						   51566 => x"0C",		-- 00c96e: 0C20            
						   51567 => x"20",
						   51568 => x"19",		-- 00c970: 1943             MOV.W   #1,R9
						   51569 => x"43",
						   51570 => x"8A",		-- 00c972: 8A93             TST.W   0x0000(R10)
						   51571 => x"93",
						   51572 => x"00",		-- 00c974: 0000            
						   51573 => x"00",
						   51574 => x"03",		-- 00c976: 0338             JL      ($C$L36)
						   51575 => x"38",
						   51576 => x"0C",		-- 00c978: 0C4A             MOV.W   R10,R12
						   51577 => x"4A",
						   51578 => x"B0",		-- 00c97a: B012             CALL    #__TI_closefile
						   51579 => x"12",
						   51580 => x"36",		-- 00c97c: 36C0            
						   51581 => x"C0",
						   51582 => x"3A",		-- 00c97e: 3A50             ADD.W   #0x000c,R10
						   51583 => x"50",
						   51584 => x"0C",		-- 00c980: 0C00            
						   51585 => x"00",
						   51586 => x"19",		-- 00c982: 1953             INC.W   R9
						   51587 => x"53",
						   51588 => x"19",		-- 00c984: 1992             CMP.W   &__TI_ft_end,R9
						   51589 => x"92",
						   51590 => x"F6",		-- 00c986: F620            
						   51591 => x"20",
						   51592 => x"F4",		-- 00c988: F43B             JL      ($C$L35)
						   51593 => x"3B",
						   51594 => x"30",		-- 00c98a: 3040             BR      #__mspabi_func_epilog_2
						   51595 => x"40",
						   51596 => x"A6",		-- 00c98c: A6CD            
						   51597 => x"CD",
						   -- Begin: finddevice
						   51598 => x"0A",		-- 00c98e: 0A12             PUSH    R10
						   51599 => x"12",
						   51600 => x"09",		-- 00c990: 0912             PUSH    R9
						   51601 => x"12",
						   51602 => x"08",		-- 00c992: 0812             PUSH    R8
						   51603 => x"12",
						   51604 => x"08",		-- 00c994: 084C             MOV.W   R12,R8
						   51605 => x"4C",
						   51606 => x"C8",		-- 00c996: C893             TST.B   0x0000(R8)
						   51607 => x"93",
						   51608 => x"00",		-- 00c998: 0000            
						   51609 => x"00",
						   51610 => x"10",		-- 00c99a: 1024             JEQ     ($C$L3)
						   51611 => x"24",
						   51612 => x"3A",		-- 00c99c: 3A40             MOV.W   #0x2092,R10
						   51613 => x"40",
						   51614 => x"92",		-- 00c99e: 9220            
						   51615 => x"20",
						   51616 => x"29",		-- 00c9a0: 2943             MOV.W   #2,R9
						   51617 => x"43",
						   51618 => x"0C",		-- 00c9a2: 0C4A             MOV.W   R10,R12
						   51619 => x"4A",
						   51620 => x"0D",		-- 00c9a4: 0D48             MOV.W   R8,R13
						   51621 => x"48",
						   51622 => x"B0",		-- 00c9a6: B012             CALL    #strcmp
						   51623 => x"12",
						   51624 => x"C2",		-- 00c9a8: C2CC            
						   51625 => x"CC",
						   51626 => x"0C",		-- 00c9aa: 0C93             TST.W   R12
						   51627 => x"93",
						   51628 => x"03",		-- 00c9ac: 0320             JNE     ($C$L2)
						   51629 => x"20",
						   51630 => x"0C",		-- 00c9ae: 0C4A             MOV.W   R10,R12
						   51631 => x"4A",
						   51632 => x"30",		-- 00c9b0: 3040             BR      #__mspabi_func_epilog_3
						   51633 => x"40",
						   51634 => x"A4",		-- 00c9b2: A4CD            
						   51635 => x"CD",
						   51636 => x"3A",		-- 00c9b4: 3A50             ADD.W   #0x001a,R10
						   51637 => x"50",
						   51638 => x"1A",		-- 00c9b6: 1A00            
						   51639 => x"00",
						   51640 => x"19",		-- 00c9b8: 1983             DEC.W   R9
						   51641 => x"83",
						   51642 => x"F3",		-- 00c9ba: F323             JNE     ($C$L1)
						   51643 => x"23",
						   51644 => x"0C",		-- 00c9bc: 0C43             CLR.W   R12
						   51645 => x"43",
						   51646 => x"30",		-- 00c9be: 3040             BR      #__mspabi_func_epilog_3
						   51647 => x"40",
						   51648 => x"A4",		-- 00c9c0: A4CD            
						   51649 => x"CD",
						   -- Begin: __TI_writemsg
						   51650 => x"82",		-- 00c9c2: 824F             MOV.W   R15,&_CIOBUF_
						   51651 => x"4F",
						   51652 => x"00",		-- 00c9c4: 0080            
						   51653 => x"80",
						   51654 => x"C2",		-- 00c9c6: C24C             MOV.B   R12,&0x8002
						   51655 => x"4C",
						   51656 => x"02",		-- 00c9c8: 0280            
						   51657 => x"80",
						   51658 => x"3C",		-- 00c9ca: 3C40             MOV.W   #0x8003,R12
						   51659 => x"40",
						   51660 => x"03",		-- 00c9cc: 0380            
						   51661 => x"80",
						   51662 => x"3B",		-- 00c9ce: 3B42             MOV.W   #8,R11
						   51663 => x"42",
						   51664 => x"1C",		-- 00c9d0: 1C53             INC.W   R12
						   51665 => x"53",
						   51666 => x"FC",		-- 00c9d2: FC4D             MOV.B   @R13+,0xffff(R12)
						   51667 => x"4D",
						   51668 => x"FF",		-- 00c9d4: FFFF            
						   51669 => x"FF",
						   51670 => x"1B",		-- 00c9d6: 1B83             DEC.W   R11
						   51671 => x"83",
						   51672 => x"FB",		-- 00c9d8: FB23             JNE     ($C$L1)
						   51673 => x"23",
						   51674 => x"0F",		-- 00c9da: 0F93             TST.W   R15
						   51675 => x"93",
						   51676 => x"07",		-- 00c9dc: 0724             JEQ     (C$$IO$$)
						   51677 => x"24",
						   51678 => x"3D",		-- 00c9de: 3D40             MOV.W   #0x800b,R13
						   51679 => x"40",
						   51680 => x"0B",		-- 00c9e0: 0B80            
						   51681 => x"80",
						   51682 => x"1D",		-- 00c9e2: 1D53             INC.W   R13
						   51683 => x"53",
						   51684 => x"FD",		-- 00c9e4: FD4E             MOV.B   @R14+,0xffff(R13)
						   51685 => x"4E",
						   51686 => x"FF",		-- 00c9e6: FFFF            
						   51687 => x"FF",
						   51688 => x"1F",		-- 00c9e8: 1F83             DEC.W   R15
						   51689 => x"83",
						   51690 => x"FB",		-- 00c9ea: FB23             JNE     ($C$L2)
						   51691 => x"23",
						   51692 => x"03",		-- 00c9ec: 0343             NOP     
						   51693 => x"43",
						   51694 => x"30",		-- 00c9ee: 3041             RET     
						   51695 => x"41",
						   -- Begin: __mspabi_subd
						   51696 => x"31",		-- 00c9f0: 3182             SUB.W   #8,SP
						   51697 => x"82",
						   51698 => x"81",		-- 00c9f2: 814C             MOV.W   R12,0x0000(SP)
						   51699 => x"4C",
						   51700 => x"00",		-- 00c9f4: 0000            
						   51701 => x"00",
						   51702 => x"81",		-- 00c9f6: 814D             MOV.W   R13,0x0002(SP)
						   51703 => x"4D",
						   51704 => x"02",		-- 00c9f8: 0200            
						   51705 => x"00",
						   51706 => x"81",		-- 00c9fa: 814E             MOV.W   R14,0x0004(SP)
						   51707 => x"4E",
						   51708 => x"04",		-- 00c9fc: 0400            
						   51709 => x"00",
						   51710 => x"81",		-- 00c9fe: 814F             MOV.W   R15,0x0006(SP)
						   51711 => x"4F",
						   51712 => x"06",		-- 00ca00: 0600            
						   51713 => x"00",
						   51714 => x"F1",		-- 00ca02: F1E0             XOR.B   #0x0080,0x0007(SP)
						   51715 => x"E0",
						   51716 => x"80",		-- 00ca04: 8000            
						   51717 => x"00",
						   51718 => x"07",		-- 00ca06: 0700            
						   51719 => x"00",
						   51720 => x"2C",		-- 00ca08: 2C41             MOV.W   @SP,R12
						   51721 => x"41",
						   51722 => x"1D",		-- 00ca0a: 1D41             MOV.W   0x0002(SP),R13
						   51723 => x"41",
						   51724 => x"02",		-- 00ca0c: 0200            
						   51725 => x"00",
						   51726 => x"1E",		-- 00ca0e: 1E41             MOV.W   0x0004(SP),R14
						   51727 => x"41",
						   51728 => x"04",		-- 00ca10: 0400            
						   51729 => x"00",
						   51730 => x"1F",		-- 00ca12: 1F41             MOV.W   0x0006(SP),R15
						   51731 => x"41",
						   51732 => x"06",		-- 00ca14: 0600            
						   51733 => x"00",
						   51734 => x"B0",		-- 00ca16: B012             CALL    #__mspabi_addd
						   51735 => x"12",
						   51736 => x"64",		-- 00ca18: 6486            
						   51737 => x"86",
						   51738 => x"31",		-- 00ca1a: 3152             ADD.W   #8,SP
						   51739 => x"52",
						   51740 => x"30",		-- 00ca1c: 3041             RET     
						   51741 => x"41",
						   -- Begin: copysignl
						   -- Begin: copysign
						   51742 => x"0A",		-- 00ca1e: 0A12             PUSH    R10
						   51743 => x"12",
						   51744 => x"1A",		-- 00ca20: 1A41             MOV.W   0x0008(SP),R10
						   51745 => x"41",
						   51746 => x"08",		-- 00ca22: 0800            
						   51747 => x"00",
						   51748 => x"1B",		-- 00ca24: 1B41             MOV.W   0x000a(SP),R11
						   51749 => x"41",
						   51750 => x"0A",		-- 00ca26: 0A00            
						   51751 => x"00",
						   51752 => x"0A",		-- 00ca28: 0AF3             AND.W   #0,R10
						   51753 => x"F3",
						   51754 => x"3B",		-- 00ca2a: 3BF0             AND.W   #0x8000,R11
						   51755 => x"F0",
						   51756 => x"00",		-- 00ca2c: 0080            
						   51757 => x"80",
						   51758 => x"3E",		-- 00ca2e: 3EF3             AND.W   #-1,R14
						   51759 => x"F3",
						   51760 => x"3F",		-- 00ca30: 3FF0             AND.W   #0x7fff,R15
						   51761 => x"F0",
						   51762 => x"FF",		-- 00ca32: FF7F            
						   51763 => x"7F",
						   51764 => x"0E",		-- 00ca34: 0EDA             BIS.W   R10,R14
						   51765 => x"DA",
						   51766 => x"0F",		-- 00ca36: 0FDB             BIS.W   R11,R15
						   51767 => x"DB",
						   51768 => x"0B",		-- 00ca38: 0B43             CLR.W   R11
						   51769 => x"43",
						   51770 => x"0B",		-- 00ca3a: 0BDD             BIS.W   R13,R11
						   51771 => x"DD",
						   51772 => x"0D",		-- 00ca3c: 0D43             CLR.W   R13
						   51773 => x"43",
						   51774 => x"0D",		-- 00ca3e: 0DDC             BIS.W   R12,R13
						   51775 => x"DC",
						   51776 => x"0E",		-- 00ca40: 0ED3             BIS.W   #0,R14
						   51777 => x"D3",
						   51778 => x"0F",		-- 00ca42: 0FD3             BIS.W   #0,R15
						   51779 => x"D3",
						   51780 => x"0C",		-- 00ca44: 0C4D             MOV.W   R13,R12
						   51781 => x"4D",
						   51782 => x"0D",		-- 00ca46: 0D4B             MOV.W   R11,R13
						   51783 => x"4B",
						   51784 => x"3A",		-- 00ca48: 3A41             POP.W   R10
						   51785 => x"41",
						   51786 => x"30",		-- 00ca4a: 3041             RET     
						   51787 => x"41",
						   -- Begin: __TI_readmsg
						   51788 => x"1F",		-- 00ca4c: 1F42             MOV.W   &_CIOBUF_,R15
						   51789 => x"42",
						   51790 => x"00",		-- 00ca4e: 0080            
						   51791 => x"80",
						   51792 => x"3B",		-- 00ca50: 3B40             MOV.W   #0x8002,R11
						   51793 => x"40",
						   51794 => x"02",		-- 00ca52: 0280            
						   51795 => x"80",
						   51796 => x"3E",		-- 00ca54: 3E42             MOV.W   #8,R14
						   51797 => x"42",
						   51798 => x"1C",		-- 00ca56: 1C53             INC.W   R12
						   51799 => x"53",
						   51800 => x"FC",		-- 00ca58: FC4B             MOV.B   @R11+,0xffff(R12)
						   51801 => x"4B",
						   51802 => x"FF",		-- 00ca5a: FFFF            
						   51803 => x"FF",
						   51804 => x"1E",		-- 00ca5c: 1E83             DEC.W   R14
						   51805 => x"83",
						   51806 => x"FB",		-- 00ca5e: FB23             JNE     ($C$L4)
						   51807 => x"23",
						   51808 => x"0D",		-- 00ca60: 0D93             TST.W   R13
						   51809 => x"93",
						   51810 => x"09",		-- 00ca62: 0924             JEQ     ($C$L6)
						   51811 => x"24",
						   51812 => x"0F",		-- 00ca64: 0F93             TST.W   R15
						   51813 => x"93",
						   51814 => x"07",		-- 00ca66: 0724             JEQ     ($C$L6)
						   51815 => x"24",
						   51816 => x"3E",		-- 00ca68: 3E40             MOV.W   #0x800a,R14
						   51817 => x"40",
						   51818 => x"0A",		-- 00ca6a: 0A80            
						   51819 => x"80",
						   51820 => x"1D",		-- 00ca6c: 1D53             INC.W   R13
						   51821 => x"53",
						   51822 => x"FD",		-- 00ca6e: FD4E             MOV.B   @R14+,0xffff(R13)
						   51823 => x"4E",
						   51824 => x"FF",		-- 00ca70: FFFF            
						   51825 => x"FF",
						   51826 => x"1F",		-- 00ca72: 1F83             DEC.W   R15
						   51827 => x"83",
						   51828 => x"FB",		-- 00ca74: FB23             JNE     ($C$L5)
						   51829 => x"23",
						   51830 => x"30",		-- 00ca76: 3041             RET     
						   51831 => x"41",
						   -- Begin: __mspabi_srai
						   51832 => x"3D",		-- 00ca78: 3DF0             AND.W   #0x000f,R13
						   51833 => x"F0",
						   51834 => x"0F",		-- 00ca7a: 0F00            
						   51835 => x"00",
						   51836 => x"3D",		-- 00ca7c: 3DE0             XOR.W   #0x000f,R13
						   51837 => x"E0",
						   51838 => x"0F",		-- 00ca7e: 0F00            
						   51839 => x"00",
						   51840 => x"0D",		-- 00ca80: 0D5D             RLA.W   R13
						   51841 => x"5D",
						   51842 => x"00",		-- 00ca82: 005D             ADD.W   R13,PC
						   51843 => x"5D",
						   -- Begin: __mspabi_srai_15
						   51844 => x"0C",		-- 00ca84: 0C11             RRA     R12
						   51845 => x"11",
						   -- Begin: __mspabi_srai_14
						   51846 => x"0C",		-- 00ca86: 0C11             RRA     R12
						   51847 => x"11",
						   -- Begin: __mspabi_srai_13
						   51848 => x"0C",		-- 00ca88: 0C11             RRA     R12
						   51849 => x"11",
						   -- Begin: __mspabi_srai_12
						   51850 => x"0C",		-- 00ca8a: 0C11             RRA     R12
						   51851 => x"11",
						   -- Begin: __mspabi_srai_11
						   51852 => x"0C",		-- 00ca8c: 0C11             RRA     R12
						   51853 => x"11",
						   -- Begin: __mspabi_srai_10
						   51854 => x"0C",		-- 00ca8e: 0C11             RRA     R12
						   51855 => x"11",
						   -- Begin: __mspabi_srai_9
						   51856 => x"0C",		-- 00ca90: 0C11             RRA     R12
						   51857 => x"11",
						   -- Begin: __mspabi_srai_8
						   51858 => x"0C",		-- 00ca92: 0C11             RRA     R12
						   51859 => x"11",
						   -- Begin: __mspabi_srai_7
						   51860 => x"0C",		-- 00ca94: 0C11             RRA     R12
						   51861 => x"11",
						   -- Begin: __mspabi_srai_6
						   51862 => x"0C",		-- 00ca96: 0C11             RRA     R12
						   51863 => x"11",
						   -- Begin: __mspabi_srai_5
						   51864 => x"0C",		-- 00ca98: 0C11             RRA     R12
						   51865 => x"11",
						   -- Begin: __mspabi_srai_4
						   51866 => x"0C",		-- 00ca9a: 0C11             RRA     R12
						   51867 => x"11",
						   -- Begin: __mspabi_srai_3
						   51868 => x"0C",		-- 00ca9c: 0C11             RRA     R12
						   51869 => x"11",
						   -- Begin: __mspabi_srai_2
						   51870 => x"0C",		-- 00ca9e: 0C11             RRA     R12
						   51871 => x"11",
						   -- Begin: __mspabi_srai_1
						   51872 => x"0C",		-- 00caa0: 0C11             RRA     R12
						   51873 => x"11",
						   51874 => x"30",		-- 00caa2: 3041             RET     
						   51875 => x"41",
						   -- Begin: __mspabi_slli
						   51876 => x"3D",		-- 00caa4: 3DF0             AND.W   #0x000f,R13
						   51877 => x"F0",
						   51878 => x"0F",		-- 00caa6: 0F00            
						   51879 => x"00",
						   51880 => x"3D",		-- 00caa8: 3DE0             XOR.W   #0x000f,R13
						   51881 => x"E0",
						   51882 => x"0F",		-- 00caaa: 0F00            
						   51883 => x"00",
						   51884 => x"0D",		-- 00caac: 0D5D             RLA.W   R13
						   51885 => x"5D",
						   51886 => x"00",		-- 00caae: 005D             ADD.W   R13,PC
						   51887 => x"5D",
						   -- Begin: __mspabi_slli_15
						   51888 => x"0C",		-- 00cab0: 0C5C             RLA.W   R12
						   51889 => x"5C",
						   -- Begin: __mspabi_slli_14
						   51890 => x"0C",		-- 00cab2: 0C5C             RLA.W   R12
						   51891 => x"5C",
						   -- Begin: __mspabi_slli_13
						   51892 => x"0C",		-- 00cab4: 0C5C             RLA.W   R12
						   51893 => x"5C",
						   -- Begin: __mspabi_slli_12
						   51894 => x"0C",		-- 00cab6: 0C5C             RLA.W   R12
						   51895 => x"5C",
						   -- Begin: __mspabi_slli_11
						   51896 => x"0C",		-- 00cab8: 0C5C             RLA.W   R12
						   51897 => x"5C",
						   -- Begin: __mspabi_slli_10
						   51898 => x"0C",		-- 00caba: 0C5C             RLA.W   R12
						   51899 => x"5C",
						   -- Begin: __mspabi_slli_9
						   51900 => x"0C",		-- 00cabc: 0C5C             RLA.W   R12
						   51901 => x"5C",
						   -- Begin: __mspabi_slli_8
						   51902 => x"0C",		-- 00cabe: 0C5C             RLA.W   R12
						   51903 => x"5C",
						   -- Begin: __mspabi_slli_7
						   51904 => x"0C",		-- 00cac0: 0C5C             RLA.W   R12
						   51905 => x"5C",
						   -- Begin: __mspabi_slli_6
						   51906 => x"0C",		-- 00cac2: 0C5C             RLA.W   R12
						   51907 => x"5C",
						   -- Begin: __mspabi_slli_5
						   51908 => x"0C",		-- 00cac4: 0C5C             RLA.W   R12
						   51909 => x"5C",
						   -- Begin: __mspabi_slli_4
						   51910 => x"0C",		-- 00cac6: 0C5C             RLA.W   R12
						   51911 => x"5C",
						   -- Begin: __mspabi_slli_3
						   51912 => x"0C",		-- 00cac8: 0C5C             RLA.W   R12
						   51913 => x"5C",
						   -- Begin: __mspabi_slli_2
						   51914 => x"0C",		-- 00caca: 0C5C             RLA.W   R12
						   51915 => x"5C",
						   -- Begin: __mspabi_slli_1
						   51916 => x"0C",		-- 00cacc: 0C5C             RLA.W   R12
						   51917 => x"5C",
						   51918 => x"30",		-- 00cace: 3041             RET     
						   51919 => x"41",
						   -- Begin: strncpy
						   51920 => x"0E",		-- 00cad0: 0E93             TST.W   R14
						   51921 => x"93",
						   51922 => x"13",		-- 00cad2: 1324             JEQ     ($C$L4)
						   51923 => x"24",
						   51924 => x"0F",		-- 00cad4: 0F4C             MOV.W   R12,R15
						   51925 => x"4C",
						   51926 => x"6B",		-- 00cad6: 6B4D             MOV.B   @R13,R11
						   51927 => x"4D",
						   51928 => x"1F",		-- 00cad8: 1F53             INC.W   R15
						   51929 => x"53",
						   51930 => x"CF",		-- 00cada: CF4B             MOV.B   R11,0xffff(R15)
						   51931 => x"4B",
						   51932 => x"FF",		-- 00cadc: FFFF            
						   51933 => x"FF",
						   51934 => x"0B",		-- 00cade: 0B93             TST.W   R11
						   51935 => x"93",
						   51936 => x"03",		-- 00cae0: 0324             JEQ     ($C$L2)
						   51937 => x"24",
						   51938 => x"1D",		-- 00cae2: 1D53             INC.W   R13
						   51939 => x"53",
						   51940 => x"1E",		-- 00cae4: 1E83             DEC.W   R14
						   51941 => x"83",
						   51942 => x"F7",		-- 00cae6: F723             JNE     ($C$L1)
						   51943 => x"23",
						   51944 => x"0D",		-- 00cae8: 0D4E             MOV.W   R14,R13
						   51945 => x"4E",
						   51946 => x"1E",		-- 00caea: 1E83             DEC.W   R14
						   51947 => x"83",
						   51948 => x"2D",		-- 00caec: 2D93             CMP.W   #2,R13
						   51949 => x"93",
						   51950 => x"05",		-- 00caee: 0528             JLO     ($C$L4)
						   51951 => x"28",
						   51952 => x"1F",		-- 00caf0: 1F53             INC.W   R15
						   51953 => x"53",
						   51954 => x"CF",		-- 00caf2: CF43             CLR.B   0xffff(R15)
						   51955 => x"43",
						   51956 => x"FF",		-- 00caf4: FFFF            
						   51957 => x"FF",
						   51958 => x"1E",		-- 00caf6: 1E83             DEC.W   R14
						   51959 => x"83",
						   51960 => x"FB",		-- 00caf8: FB23             JNE     ($C$L3)
						   51961 => x"23",
						   51962 => x"30",		-- 00cafa: 3041             RET     
						   51963 => x"41",
						   -- Begin: __mspabi_negd
						   51964 => x"31",		-- 00cafc: 3182             SUB.W   #8,SP
						   51965 => x"82",
						   51966 => x"81",		-- 00cafe: 814C             MOV.W   R12,0x0000(SP)
						   51967 => x"4C",
						   51968 => x"00",		-- 00cb00: 0000            
						   51969 => x"00",
						   51970 => x"81",		-- 00cb02: 814D             MOV.W   R13,0x0002(SP)
						   51971 => x"4D",
						   51972 => x"02",		-- 00cb04: 0200            
						   51973 => x"00",
						   51974 => x"81",		-- 00cb06: 814E             MOV.W   R14,0x0004(SP)
						   51975 => x"4E",
						   51976 => x"04",		-- 00cb08: 0400            
						   51977 => x"00",
						   51978 => x"81",		-- 00cb0a: 814F             MOV.W   R15,0x0006(SP)
						   51979 => x"4F",
						   51980 => x"06",		-- 00cb0c: 0600            
						   51981 => x"00",
						   51982 => x"F1",		-- 00cb0e: F1E0             XOR.B   #0x0080,0x0007(SP)
						   51983 => x"E0",
						   51984 => x"80",		-- 00cb10: 8000            
						   51985 => x"00",
						   51986 => x"07",		-- 00cb12: 0700            
						   51987 => x"00",
						   51988 => x"2C",		-- 00cb14: 2C41             MOV.W   @SP,R12
						   51989 => x"41",
						   51990 => x"1D",		-- 00cb16: 1D41             MOV.W   0x0002(SP),R13
						   51991 => x"41",
						   51992 => x"02",		-- 00cb18: 0200            
						   51993 => x"00",
						   51994 => x"1E",		-- 00cb1a: 1E41             MOV.W   0x0004(SP),R14
						   51995 => x"41",
						   51996 => x"04",		-- 00cb1c: 0400            
						   51997 => x"00",
						   51998 => x"1F",		-- 00cb1e: 1F41             MOV.W   0x0006(SP),R15
						   51999 => x"41",
						   52000 => x"06",		-- 00cb20: 0600            
						   52001 => x"00",
						   52002 => x"31",		-- 00cb22: 3152             ADD.W   #8,SP
						   52003 => x"52",
						   52004 => x"30",		-- 00cb24: 3041             RET     
						   52005 => x"41",
						   -- Begin: __mspabi_fixdi
						   52006 => x"B0",		-- 00cb26: B012             CALL    #__mspabi_fixdli
						   52007 => x"12",
						   52008 => x"A8",		-- 00cb28: A8C0            
						   52009 => x"C0",
						   52010 => x"0D",		-- 00cb2a: 0D93             TST.W   R13
						   52011 => x"93",
						   52012 => x"07",		-- 00cb2c: 0738             JL      ($C$L7)
						   52013 => x"38",
						   52014 => x"03",		-- 00cb2e: 0320             JNE     ($C$L6)
						   52015 => x"20",
						   52016 => x"3C",		-- 00cb30: 3C90             CMP.W   #0x8000,R12
						   52017 => x"90",
						   52018 => x"00",		-- 00cb32: 0080            
						   52019 => x"80",
						   52020 => x"03",		-- 00cb34: 0328             JLO     ($C$L7)
						   52021 => x"28",
						   52022 => x"3C",		-- 00cb36: 3C40             MOV.W   #0x7fff,R12
						   52023 => x"40",
						   52024 => x"FF",		-- 00cb38: FF7F            
						   52025 => x"7F",
						   52026 => x"30",		-- 00cb3a: 3041             RET     
						   52027 => x"41",
						   52028 => x"3D",		-- 00cb3c: 3D93             CMP.W   #-1,R13
						   52029 => x"93",
						   52030 => x"04",		-- 00cb3e: 0438             JL      ($C$L8)
						   52031 => x"38",
						   52032 => x"05",		-- 00cb40: 0520             JNE     ($C$L9)
						   52033 => x"20",
						   52034 => x"3C",		-- 00cb42: 3C90             CMP.W   #0x8000,R12
						   52035 => x"90",
						   52036 => x"00",		-- 00cb44: 0080            
						   52037 => x"80",
						   52038 => x"02",		-- 00cb46: 022C             JHS     ($C$L9)
						   52039 => x"2C",
						   52040 => x"3C",		-- 00cb48: 3C40             MOV.W   #0x8000,R12
						   52041 => x"40",
						   52042 => x"00",		-- 00cb4a: 0080            
						   52043 => x"80",
						   52044 => x"30",		-- 00cb4c: 3041             RET     
						   52045 => x"41",
						   -- Begin: free_list_insert
						   52046 => x"2F",		-- 00cb4e: 2F4C             MOV.W   @R12,R15
						   52047 => x"4C",
						   52048 => x"1F",		-- 00cb50: 1FC3             BIC.W   #1,R15
						   52049 => x"C3",
						   52050 => x"3E",		-- 00cb52: 3E40             MOV.W   #0x21a6,R14
						   52051 => x"40",
						   52052 => x"A6",		-- 00cb54: A621            
						   52053 => x"21",
						   52054 => x"03",		-- 00cb56: 033C             JMP     ($C$L5)
						   52055 => x"3C",
						   52056 => x"2D",		-- 00cb58: 2D42             MOV.W   #4,R13
						   52057 => x"42",
						   52058 => x"2D",		-- 00cb5a: 2D5E             ADD.W   @R14,R13
						   52059 => x"5E",
						   52060 => x"0E",		-- 00cb5c: 0E4D             MOV.W   R13,R14
						   52061 => x"4D",
						   52062 => x"2D",		-- 00cb5e: 2D4E             MOV.W   @R14,R13
						   52063 => x"4E",
						   52064 => x"0D",		-- 00cb60: 0D93             TST.W   R13
						   52065 => x"93",
						   52066 => x"04",		-- 00cb62: 0424             JEQ     ($C$L6)
						   52067 => x"24",
						   52068 => x"2D",		-- 00cb64: 2D4D             MOV.W   @R13,R13
						   52069 => x"4D",
						   52070 => x"1D",		-- 00cb66: 1DC3             BIC.W   #1,R13
						   52071 => x"C3",
						   52072 => x"0D",		-- 00cb68: 0D9F             CMP.W   R15,R13
						   52073 => x"9F",
						   52074 => x"F6",		-- 00cb6a: F62B             JLO     ($C$L4)
						   52075 => x"2B",
						   52076 => x"AC",		-- 00cb6c: AC4E             MOV.W   @R14,0x0004(R12)
						   52077 => x"4E",
						   52078 => x"04",		-- 00cb6e: 0400            
						   52079 => x"00",
						   52080 => x"8E",		-- 00cb70: 8E4C             MOV.W   R12,0x0000(R14)
						   52081 => x"4C",
						   52082 => x"00",		-- 00cb72: 0000            
						   52083 => x"00",
						   52084 => x"30",		-- 00cb74: 3041             RET     
						   52085 => x"41",
						   -- Begin: remove
						   -- Begin: unlink
						   52086 => x"0A",		-- 00cb76: 0A12             PUSH    R10
						   52087 => x"12",
						   52088 => x"21",		-- 00cb78: 2183             DECD.W  SP
						   52089 => x"83",
						   52090 => x"81",		-- 00cb7a: 814C             MOV.W   R12,0x0000(SP)
						   52091 => x"4C",
						   52092 => x"00",		-- 00cb7c: 0000            
						   52093 => x"00",
						   52094 => x"92",		-- 00cb7e: 9212             CALL    &_lock
						   52095 => x"12",
						   52096 => x"F2",		-- 00cb80: F220            
						   52097 => x"20",
						   52098 => x"0C",		-- 00cb82: 0C41             MOV.W   SP,R12
						   52099 => x"41",
						   52100 => x"B0",		-- 00cb84: B012             CALL    #getdevice
						   52101 => x"12",
						   52102 => x"9E",		-- 00cb86: 9EC4            
						   52103 => x"C4",
						   52104 => x"0F",		-- 00cb88: 0F4C             MOV.W   R12,R15
						   52105 => x"4C",
						   52106 => x"2C",		-- 00cb8a: 2C41             MOV.W   @SP,R12
						   52107 => x"41",
						   52108 => x"9F",		-- 00cb8c: 9F12             CALL    0x0016(R15)
						   52109 => x"12",
						   52110 => x"16",		-- 00cb8e: 1600            
						   52111 => x"00",
						   52112 => x"0A",		-- 00cb90: 0A4C             MOV.W   R12,R10
						   52113 => x"4C",
						   52114 => x"92",		-- 00cb92: 9212             CALL    &_unlock
						   52115 => x"12",
						   52116 => x"F4",		-- 00cb94: F420            
						   52117 => x"20",
						   52118 => x"0C",		-- 00cb96: 0C4A             MOV.W   R10,R12
						   52119 => x"4A",
						   52120 => x"21",		-- 00cb98: 2153             INCD.W  SP
						   52121 => x"53",
						   52122 => x"3A",		-- 00cb9a: 3A41             POP.W   R10
						   52123 => x"41",
						   52124 => x"30",		-- 00cb9c: 3041             RET     
						   52125 => x"41",
						   -- Begin: lseek
						   52126 => x"0C",		-- 00cb9e: 0C93             TST.W   R12
						   52127 => x"93",
						   52128 => x"0E",		-- 00cba0: 0E38             JL      ($C$L1)
						   52129 => x"38",
						   52130 => x"3C",		-- 00cba2: 3C90             CMP.W   #0x000a,R12
						   52131 => x"90",
						   52132 => x"0A",		-- 00cba4: 0A00            
						   52133 => x"00",
						   52134 => x"0B",		-- 00cba6: 0B34             JGE     ($C$L1)
						   52135 => x"34",
						   52136 => x"0C",		-- 00cba8: 0C5C             RLA.W   R12
						   52137 => x"5C",
						   52138 => x"0C",		-- 00cbaa: 0C5C             RLA.W   R12
						   52139 => x"5C",
						   52140 => x"3C",		-- 00cbac: 3C50             ADD.W   #0x20c6,R12
						   52141 => x"50",
						   52142 => x"C6",		-- 00cbae: C620            
						   52143 => x"20",
						   52144 => x"2B",		-- 00cbb0: 2B4C             MOV.W   @R12,R11
						   52145 => x"4C",
						   52146 => x"0B",		-- 00cbb2: 0B93             TST.W   R11
						   52147 => x"93",
						   52148 => x"04",		-- 00cbb4: 0424             JEQ     ($C$L1)
						   52149 => x"24",
						   52150 => x"1C",		-- 00cbb6: 1C4C             MOV.W   0x0002(R12),R12
						   52151 => x"4C",
						   52152 => x"02",		-- 00cbb8: 0200            
						   52153 => x"00",
						   52154 => x"10",		-- 00cbba: 104B             BR      0x0014(R11)
						   52155 => x"4B",
						   52156 => x"14",		-- 00cbbc: 1400            
						   52157 => x"00",
						   52158 => x"3C",		-- 00cbbe: 3C43             MOV.W   #-1,R12
						   52159 => x"43",
						   52160 => x"3D",		-- 00cbc0: 3D43             MOV.W   #-1,R13
						   52161 => x"43",
						   52162 => x"30",		-- 00cbc2: 3041             RET     
						   52163 => x"41",
						   -- Begin: __mspabi_mpyl
						   -- Begin: __mspabi_mpyl_sw
						   52164 => x"0A",		-- 00cbc4: 0A12             PUSH    R10
						   52165 => x"12",
						   52166 => x"0A",		-- 00cbc6: 0A43             CLR.W   R10
						   52167 => x"43",
						   52168 => x"0B",		-- 00cbc8: 0B43             CLR.W   R11
						   52169 => x"43",
						   -- Begin: mpyl_add_loop
						   52170 => x"12",		-- 00cbca: 12C3             CLRC    
						   52171 => x"C3",
						   52172 => x"0D",		-- 00cbcc: 0D10             RRC     R13
						   52173 => x"10",
						   52174 => x"0C",		-- 00cbce: 0C10             RRC     R12
						   52175 => x"10",
						   52176 => x"02",		-- 00cbd0: 0228             JLO     (shift_test_mpyl)
						   52177 => x"28",
						   52178 => x"0A",		-- 00cbd2: 0A5E             ADD.W   R14,R10
						   52179 => x"5E",
						   52180 => x"0B",		-- 00cbd4: 0B6F             ADDC.W  R15,R11
						   52181 => x"6F",
						   -- Begin: shift_test_mpyl
						   52182 => x"0E",		-- 00cbd6: 0E5E             RLA.W   R14
						   52183 => x"5E",
						   52184 => x"0F",		-- 00cbd8: 0F6F             RLC.W   R15
						   52185 => x"6F",
						   52186 => x"0D",		-- 00cbda: 0D93             TST.W   R13
						   52187 => x"93",
						   52188 => x"F6",		-- 00cbdc: F623             JNE     (mpyl_add_loop)
						   52189 => x"23",
						   52190 => x"0C",		-- 00cbde: 0C93             TST.W   R12
						   52191 => x"93",
						   52192 => x"F4",		-- 00cbe0: F423             JNE     (mpyl_add_loop)
						   52193 => x"23",
						   52194 => x"0C",		-- 00cbe2: 0C4A             MOV.W   R10,R12
						   52195 => x"4A",
						   52196 => x"0D",		-- 00cbe4: 0D4B             MOV.W   R11,R13
						   52197 => x"4B",
						   52198 => x"3A",		-- 00cbe6: 3A41             POP.W   R10
						   52199 => x"41",
						   52200 => x"30",		-- 00cbe8: 3041             RET     
						   52201 => x"41",
						   -- Begin: write
						   52202 => x"0C",		-- 00cbea: 0C93             TST.W   R12
						   52203 => x"93",
						   52204 => x"0E",		-- 00cbec: 0E38             JL      ($C$L1)
						   52205 => x"38",
						   52206 => x"3C",		-- 00cbee: 3C90             CMP.W   #0x000a,R12
						   52207 => x"90",
						   52208 => x"0A",		-- 00cbf0: 0A00            
						   52209 => x"00",
						   52210 => x"0B",		-- 00cbf2: 0B34             JGE     ($C$L1)
						   52211 => x"34",
						   52212 => x"0C",		-- 00cbf4: 0C5C             RLA.W   R12
						   52213 => x"5C",
						   52214 => x"0C",		-- 00cbf6: 0C5C             RLA.W   R12
						   52215 => x"5C",
						   52216 => x"3C",		-- 00cbf8: 3C50             ADD.W   #0x20c6,R12
						   52217 => x"50",
						   52218 => x"C6",		-- 00cbfa: C620            
						   52219 => x"20",
						   52220 => x"2F",		-- 00cbfc: 2F4C             MOV.W   @R12,R15
						   52221 => x"4C",
						   52222 => x"0F",		-- 00cbfe: 0F93             TST.W   R15
						   52223 => x"93",
						   52224 => x"04",		-- 00cc00: 0424             JEQ     ($C$L1)
						   52225 => x"24",
						   52226 => x"1C",		-- 00cc02: 1C4C             MOV.W   0x0002(R12),R12
						   52227 => x"4C",
						   52228 => x"02",		-- 00cc04: 0200            
						   52229 => x"00",
						   52230 => x"10",		-- 00cc06: 104F             BR      0x0012(R15)
						   52231 => x"4F",
						   52232 => x"12",		-- 00cc08: 1200            
						   52233 => x"00",
						   52234 => x"3C",		-- 00cc0a: 3C43             MOV.W   #-1,R12
						   52235 => x"43",
						   52236 => x"30",		-- 00cc0c: 3041             RET     
						   52237 => x"41",
						   -- Begin: __mspabi_mpyul
						   -- Begin: __mspabi_mpyul_sw
						   52238 => x"0B",		-- 00cc0e: 0B4C             MOV.W   R12,R11
						   52239 => x"4C",
						   52240 => x"0E",		-- 00cc10: 0E4D             MOV.W   R13,R14
						   52241 => x"4D",
						   52242 => x"0F",		-- 00cc12: 0F43             CLR.W   R15
						   52243 => x"43",
						   52244 => x"0C",		-- 00cc14: 0C43             CLR.W   R12
						   52245 => x"43",
						   52246 => x"0D",		-- 00cc16: 0D43             CLR.W   R13
						   52247 => x"43",
						   52248 => x"12",		-- 00cc18: 12C3             CLRC    
						   52249 => x"C3",
						   52250 => x"0B",		-- 00cc1a: 0B10             RRC     R11
						   52251 => x"10",
						   52252 => x"01",		-- 00cc1c: 013C             JMP     (mpyul_add_loop1)
						   52253 => x"3C",
						   -- Begin: mpyul_add_loop
						   52254 => x"0B",		-- 00cc1e: 0B11             RRA     R11
						   52255 => x"11",
						   -- Begin: mpyul_add_loop1
						   52256 => x"02",		-- 00cc20: 0228             JLO     (shift_test_mpyul)
						   52257 => x"28",
						   52258 => x"0C",		-- 00cc22: 0C5E             ADD.W   R14,R12
						   52259 => x"5E",
						   52260 => x"0D",		-- 00cc24: 0D6F             ADDC.W  R15,R13
						   52261 => x"6F",
						   -- Begin: shift_test_mpyul
						   52262 => x"0E",		-- 00cc26: 0E5E             RLA.W   R14
						   52263 => x"5E",
						   52264 => x"0F",		-- 00cc28: 0F6F             RLC.W   R15
						   52265 => x"6F",
						   52266 => x"0B",		-- 00cc2a: 0B93             TST.W   R11
						   52267 => x"93",
						   52268 => x"F8",		-- 00cc2c: F823             JNE     (mpyul_add_loop)
						   52269 => x"23",
						   52270 => x"30",		-- 00cc2e: 3041             RET     
						   52271 => x"41",
						   -- Begin: memccpy
						   52272 => x"0A",		-- 00cc30: 0A12             PUSH    R10
						   52273 => x"12",
						   52274 => x"0F",		-- 00cc32: 0F93             TST.W   R15
						   52275 => x"93",
						   52276 => x"0B",		-- 00cc34: 0B24             JEQ     ($C$L2)
						   52277 => x"24",
						   52278 => x"4E",		-- 00cc36: 4E4E             MOV.B   R14,R14
						   52279 => x"4E",
						   52280 => x"6B",		-- 00cc38: 6B4D             MOV.B   @R13,R11
						   52281 => x"4D",
						   52282 => x"1C",		-- 00cc3a: 1C53             INC.W   R12
						   52283 => x"53",
						   52284 => x"CC",		-- 00cc3c: CC4B             MOV.B   R11,0xffff(R12)
						   52285 => x"4B",
						   52286 => x"FF",		-- 00cc3e: FFFF            
						   52287 => x"FF",
						   52288 => x"4A",		-- 00cc40: 4A4E             MOV.B   R14,R10
						   52289 => x"4E",
						   52290 => x"0B",		-- 00cc42: 0B9A             CMP.W   R10,R11
						   52291 => x"9A",
						   52292 => x"04",		-- 00cc44: 0424             JEQ     ($C$L3)
						   52293 => x"24",
						   52294 => x"1D",		-- 00cc46: 1D53             INC.W   R13
						   52295 => x"53",
						   52296 => x"1F",		-- 00cc48: 1F83             DEC.W   R15
						   52297 => x"83",
						   52298 => x"F6",		-- 00cc4a: F623             JNE     ($C$L1)
						   52299 => x"23",
						   52300 => x"0C",		-- 00cc4c: 0C43             CLR.W   R12
						   52301 => x"43",
						   52302 => x"3A",		-- 00cc4e: 3A41             POP.W   R10
						   52303 => x"41",
						   52304 => x"30",		-- 00cc50: 3041             RET     
						   52305 => x"41",
						   -- Begin: __mspabi_mpyull
						   -- Begin: __mspabi_mpyull_sw
						   52306 => x"0A",		-- 00cc52: 0A12             PUSH    R10
						   52307 => x"12",
						   52308 => x"09",		-- 00cc54: 0912             PUSH    R9
						   52309 => x"12",
						   52310 => x"08",		-- 00cc56: 0812             PUSH    R8
						   52311 => x"12",
						   52312 => x"08",		-- 00cc58: 084C             MOV.W   R12,R8
						   52313 => x"4C",
						   52314 => x"09",		-- 00cc5a: 094D             MOV.W   R13,R9
						   52315 => x"4D",
						   52316 => x"0A",		-- 00cc5c: 0A43             CLR.W   R10
						   52317 => x"43",
						   52318 => x"0B",		-- 00cc5e: 0B43             CLR.W   R11
						   52319 => x"43",
						   52320 => x"0C",		-- 00cc60: 0C4E             MOV.W   R14,R12
						   52321 => x"4E",
						   52322 => x"0D",		-- 00cc62: 0D4F             MOV.W   R15,R13
						   52323 => x"4F",
						   52324 => x"0E",		-- 00cc64: 0E43             CLR.W   R14
						   52325 => x"43",
						   52326 => x"0F",		-- 00cc66: 0F43             CLR.W   R15
						   52327 => x"43",
						   52328 => x"B0",		-- 00cc68: B012             CALL    #__mspabi_mpyll_sw
						   52329 => x"12",
						   52330 => x"F4",		-- 00cc6a: F4B1            
						   52331 => x"B1",
						   52332 => x"30",		-- 00cc6c: 3040             BR      #__mspabi_func_epilog_3
						   52333 => x"40",
						   52334 => x"A4",		-- 00cc6e: A4CD            
						   52335 => x"CD",
						   -- Begin: _c_int00_noargs
						   52336 => x"31",		-- 00cc70: 3140             MOV.W   #0x3000,SP
						   52337 => x"40",
						   52338 => x"00",		-- 00cc72: 0030            
						   52339 => x"30",
						   52340 => x"B0",		-- 00cc74: B012             CALL    #_system_pre_init
						   52341 => x"12",
						   52342 => x"04",		-- 00cc76: 04CE            
						   52343 => x"CE",
						   52344 => x"0C",		-- 00cc78: 0C93             TST.W   R12
						   52345 => x"93",
						   52346 => x"02",		-- 00cc7a: 0224             JEQ     ($C$L2)
						   52347 => x"24",
						   52348 => x"B0",		-- 00cc7c: B012             CALL    #__TI_auto_init_nobinit_nopinit
						   52349 => x"12",
						   52350 => x"E0",		-- 00cc7e: E0C7            
						   52351 => x"C7",
						   52352 => x"0C",		-- 00cc80: 0C43             CLR.W   R12
						   52353 => x"43",
						   52354 => x"B0",		-- 00cc82: B012             CALL    #main
						   52355 => x"12",
						   52356 => x"42",		-- 00cc84: 42C4            
						   52357 => x"C4",
						   52358 => x"1C",		-- 00cc86: 1C43             MOV.W   #1,R12
						   52359 => x"43",
						   52360 => x"B0",		-- 00cc88: B012             CALL    #exit
						   52361 => x"12",
						   52362 => x"9C",		-- 00cc8a: 9CC7            
						   52363 => x"C7",
						   -- Begin: free_list_remove
						   52364 => x"3F",		-- 00cc8c: 3F40             MOV.W   #0x21a6,R15
						   52365 => x"40",
						   52366 => x"A6",		-- 00cc8e: A621            
						   52367 => x"21",
						   52368 => x"02",		-- 00cc90: 023C             JMP     ($C$L2)
						   52369 => x"3C",
						   52370 => x"2F",		-- 00cc92: 2F42             MOV.W   #4,R15
						   52371 => x"42",
						   52372 => x"0F",		-- 00cc94: 0F5E             ADD.W   R14,R15
						   52373 => x"5E",
						   52374 => x"2E",		-- 00cc96: 2E4F             MOV.W   @R15,R14
						   52375 => x"4F",
						   52376 => x"0E",		-- 00cc98: 0E93             TST.W   R14
						   52377 => x"93",
						   52378 => x"05",		-- 00cc9a: 0524             JEQ     ($C$L3)
						   52379 => x"24",
						   52380 => x"0E",		-- 00cc9c: 0E9C             CMP.W   R12,R14
						   52381 => x"9C",
						   52382 => x"F9",		-- 00cc9e: F923             JNE     ($C$L1)
						   52383 => x"23",
						   52384 => x"9F",		-- 00cca0: 9F4C             MOV.W   0x0004(R12),0x0000(R15)
						   52385 => x"4C",
						   52386 => x"04",		-- 00cca2: 0400            
						   52387 => x"00",
						   52388 => x"00",		-- 00cca4: 0000            
						   52389 => x"00",
						   52390 => x"30",		-- 00cca6: 3041             RET     
						   52391 => x"41",
						   -- Begin: strchr
						   52392 => x"6F",		-- 00cca8: 6F4C             MOV.B   @R12,R15
						   52393 => x"4C",
						   52394 => x"4D",		-- 00ccaa: 4D4D             MOV.B   R13,R13
						   52395 => x"4D",
						   52396 => x"06",		-- 00ccac: 063C             JMP     ($C$L3)
						   52397 => x"3C",
						   52398 => x"0F",		-- 00ccae: 0F93             TST.W   R15
						   52399 => x"93",
						   52400 => x"02",		-- 00ccb0: 0220             JNE     ($C$L2)
						   52401 => x"20",
						   52402 => x"0C",		-- 00ccb2: 0C43             CLR.W   R12
						   52403 => x"43",
						   52404 => x"30",		-- 00ccb4: 3041             RET     
						   52405 => x"41",
						   52406 => x"1C",		-- 00ccb6: 1C53             INC.W   R12
						   52407 => x"53",
						   52408 => x"6F",		-- 00ccb8: 6F4C             MOV.B   @R12,R15
						   52409 => x"4C",
						   52410 => x"4E",		-- 00ccba: 4E4D             MOV.B   R13,R14
						   52411 => x"4D",
						   52412 => x"0F",		-- 00ccbc: 0F9E             CMP.W   R14,R15
						   52413 => x"9E",
						   52414 => x"F7",		-- 00ccbe: F723             JNE     ($C$L1)
						   52415 => x"23",
						   52416 => x"30",		-- 00ccc0: 3041             RET     
						   52417 => x"41",
						   -- Begin: strcmp
						   52418 => x"0F",		-- 00ccc2: 0F4C             MOV.W   R12,R15
						   52419 => x"4C",
						   52420 => x"6E",		-- 00ccc4: 6E4F             MOV.B   @R15,R14
						   52421 => x"4F",
						   52422 => x"6B",		-- 00ccc6: 6B4D             MOV.B   @R13,R11
						   52423 => x"4D",
						   52424 => x"4C",		-- 00ccc8: 4C4E             MOV.B   R14,R12
						   52425 => x"4E",
						   52426 => x"0C",		-- 00ccca: 0C8B             SUB.W   R11,R12
						   52427 => x"8B",
						   52428 => x"4E",		-- 00cccc: 4E93             TST.B   R14
						   52429 => x"93",
						   52430 => x"04",		-- 00ccce: 0424             JEQ     ($C$L2)
						   52431 => x"24",
						   52432 => x"1D",		-- 00ccd0: 1D53             INC.W   R13
						   52433 => x"53",
						   52434 => x"1F",		-- 00ccd2: 1F53             INC.W   R15
						   52435 => x"53",
						   52436 => x"0C",		-- 00ccd4: 0C93             TST.W   R12
						   52437 => x"93",
						   52438 => x"F6",		-- 00ccd6: F627             JEQ     ($C$L1)
						   52439 => x"27",
						   52440 => x"30",		-- 00ccd8: 3041             RET     
						   52441 => x"41",
						   -- Begin: __mspabi_divu
						   -- Begin: __mspabi_remu
						   52442 => x"0E",		-- 00ccda: 0E43             CLR.W   R14
						   52443 => x"43",
						   52444 => x"0F",		-- 00ccdc: 0F4C             MOV.W   R12,R15
						   52445 => x"4C",
						   52446 => x"1C",		-- 00ccde: 1C43             MOV.W   #1,R12
						   52447 => x"43",
						   -- Begin: div_loop
						   52448 => x"0F",		-- 00cce0: 0F5F             RLA.W   R15
						   52449 => x"5F",
						   52450 => x"0E",		-- 00cce2: 0E6E             RLC.W   R14
						   52451 => x"6E",
						   52452 => x"0E",		-- 00cce4: 0E9D             CMP.W   R13,R14
						   52453 => x"9D",
						   52454 => x"01",		-- 00cce6: 0128             JLO     (set_quotient_bit)
						   52455 => x"28",
						   52456 => x"0E",		-- 00cce8: 0E8D             SUB.W   R13,R14
						   52457 => x"8D",
						   -- Begin: set_quotient_bit
						   52458 => x"0C",		-- 00ccea: 0C6C             RLC.W   R12
						   52459 => x"6C",
						   52460 => x"F9",		-- 00ccec: F92B             JLO     (div_loop)
						   52461 => x"2B",
						   52462 => x"30",		-- 00ccee: 3041             RET     
						   52463 => x"41",
						   -- Begin: __TI_zero_init_nomemset
						   52464 => x"1F",		-- 00ccf0: 1F4C             MOV.W   0x0001(R12),R15
						   52465 => x"4C",
						   52466 => x"01",		-- 00ccf2: 0100            
						   52467 => x"00",
						   52468 => x"0F",		-- 00ccf4: 0F93             TST.W   R15
						   52469 => x"93",
						   52470 => x"05",		-- 00ccf6: 0524             JEQ     ($C$L2)
						   52471 => x"24",
						   52472 => x"1D",		-- 00ccf8: 1D53             INC.W   R13
						   52473 => x"53",
						   52474 => x"CD",		-- 00ccfa: CD43             CLR.B   0xffff(R13)
						   52475 => x"43",
						   52476 => x"FF",		-- 00ccfc: FFFF            
						   52477 => x"FF",
						   52478 => x"1F",		-- 00ccfe: 1F83             DEC.W   R15
						   52479 => x"83",
						   52480 => x"FB",		-- 00cd00: FB23             JNE     ($C$L1)
						   52481 => x"23",
						   52482 => x"30",		-- 00cd02: 3041             RET     
						   52483 => x"41",
						   -- Begin: memchr
						   52484 => x"0E",		-- 00cd04: 0E93             TST.W   R14
						   52485 => x"93",
						   52486 => x"06",		-- 00cd06: 0624             JEQ     ($C$L2)
						   52487 => x"24",
						   52488 => x"4D",		-- 00cd08: 4D4D             MOV.B   R13,R13
						   52489 => x"4D",
						   52490 => x"6D",		-- 00cd0a: 6D9C             CMP.B   @R12,R13
						   52491 => x"9C",
						   52492 => x"04",		-- 00cd0c: 0424             JEQ     ($C$L3)
						   52493 => x"24",
						   52494 => x"1C",		-- 00cd0e: 1C53             INC.W   R12
						   52495 => x"53",
						   52496 => x"1E",		-- 00cd10: 1E83             DEC.W   R14
						   52497 => x"83",
						   52498 => x"FB",		-- 00cd12: FB23             JNE     ($C$L1)
						   52499 => x"23",
						   52500 => x"0C",		-- 00cd14: 0C43             CLR.W   R12
						   52501 => x"43",
						   52502 => x"30",		-- 00cd16: 3041             RET     
						   52503 => x"41",
						   -- Begin: memset
						   52504 => x"0F",		-- 00cd18: 0F4C             MOV.W   R12,R15
						   52505 => x"4C",
						   52506 => x"0E",		-- 00cd1a: 0E93             TST.W   R14
						   52507 => x"93",
						   52508 => x"06",		-- 00cd1c: 0624             JEQ     ($C$L2)
						   52509 => x"24",
						   52510 => x"4D",		-- 00cd1e: 4D4D             MOV.B   R13,R13
						   52511 => x"4D",
						   52512 => x"1F",		-- 00cd20: 1F53             INC.W   R15
						   52513 => x"53",
						   52514 => x"CF",		-- 00cd22: CF4D             MOV.B   R13,0xffff(R15)
						   52515 => x"4D",
						   52516 => x"FF",		-- 00cd24: FFFF            
						   52517 => x"FF",
						   52518 => x"1E",		-- 00cd26: 1E83             DEC.W   R14
						   52519 => x"83",
						   52520 => x"FB",		-- 00cd28: FB23             JNE     ($C$L1)
						   52521 => x"23",
						   52522 => x"30",		-- 00cd2a: 3041             RET     
						   52523 => x"41",
						   -- Begin: __mspabi_mpyi
						   -- Begin: __mspabi_mpyi_sw
						   52524 => x"0E",		-- 00cd2c: 0E43             CLR.W   R14
						   52525 => x"43",
						   -- Begin: mpyi_add_loop
						   52526 => x"12",		-- 00cd2e: 12C3             CLRC    
						   52527 => x"C3",
						   52528 => x"0C",		-- 00cd30: 0C10             RRC     R12
						   52529 => x"10",
						   52530 => x"01",		-- 00cd32: 0128             JLO     (shift_test_mpyi)
						   52531 => x"28",
						   52532 => x"0E",		-- 00cd34: 0E5D             ADD.W   R13,R14
						   52533 => x"5D",
						   -- Begin: shift_test_mpyi
						   52534 => x"0D",		-- 00cd36: 0D5D             RLA.W   R13
						   52535 => x"5D",
						   52536 => x"0C",		-- 00cd38: 0C93             TST.W   R12
						   52537 => x"93",
						   52538 => x"F9",		-- 00cd3a: F923             JNE     (mpyi_add_loop)
						   52539 => x"23",
						   52540 => x"0C",		-- 00cd3c: 0C4E             MOV.W   R14,R12
						   52541 => x"4E",
						   52542 => x"30",		-- 00cd3e: 3041             RET     
						   52543 => x"41",
						   -- Begin: wcslen
						   52544 => x"0F",		-- 00cd40: 0F4C             MOV.W   R12,R15
						   52545 => x"4C",
						   52546 => x"01",		-- 00cd42: 013C             JMP     ($C$L2)
						   52547 => x"3C",
						   52548 => x"2F",		-- 00cd44: 2F53             INCD.W  R15
						   52549 => x"53",
						   52550 => x"8F",		-- 00cd46: 8F93             TST.W   0x0000(R15)
						   52551 => x"93",
						   52552 => x"00",		-- 00cd48: 0000            
						   52553 => x"00",
						   52554 => x"FC",		-- 00cd4a: FC23             JNE     ($C$L1)
						   52555 => x"23",
						   52556 => x"0F",		-- 00cd4c: 0F8C             SUB.W   R12,R15
						   52557 => x"8C",
						   52558 => x"0F",		-- 00cd4e: 0F11             RRA     R15
						   52559 => x"11",
						   52560 => x"0C",		-- 00cd50: 0C4F             MOV.W   R15,R12
						   52561 => x"4F",
						   52562 => x"30",		-- 00cd52: 3041             RET     
						   52563 => x"41",
						   -- Begin: buff_value
						   52564 => x"21",		-- 00cd54: 2183             DECD.W  SP
						   52565 => x"83",
						   52566 => x"81",		-- 00cd56: 814C             MOV.W   R12,0x0000(SP)
						   52567 => x"4C",
						   52568 => x"00",		-- 00cd58: 0000            
						   52569 => x"00",
						   52570 => x"3D",		-- 00cd5a: 3D40             MOV.W   #0x863c,R13
						   52571 => x"40",
						   52572 => x"3C",		-- 00cd5c: 3C86            
						   52573 => x"86",
						   52574 => x"B0",		-- 00cd5e: B012             CALL    #strcpy
						   52575 => x"12",
						   52576 => x"AC",		-- 00cd60: ACCD            
						   52577 => x"CD",
						   52578 => x"21",		-- 00cd62: 2153             INCD.W  SP
						   52579 => x"53",
						   52580 => x"30",		-- 00cd64: 3041             RET     
						   52581 => x"41",
						   -- Begin: __TI_decompress_none
						   52582 => x"0F",		-- 00cd66: 0F4C             MOV.W   R12,R15
						   52583 => x"4C",
						   52584 => x"0C",		-- 00cd68: 0C4D             MOV.W   R13,R12
						   52585 => x"4D",
						   52586 => x"3D",		-- 00cd6a: 3D40             MOV.W   #0x0003,R13
						   52587 => x"40",
						   52588 => x"03",		-- 00cd6c: 0300            
						   52589 => x"00",
						   52590 => x"0D",		-- 00cd6e: 0D5F             ADD.W   R15,R13
						   52591 => x"5F",
						   52592 => x"1E",		-- 00cd70: 1E4F             MOV.W   0x0001(R15),R14
						   52593 => x"4F",
						   52594 => x"01",		-- 00cd72: 0100            
						   52595 => x"00",
						   52596 => x"30",		-- 00cd74: 3040             BR      #memcpy
						   52597 => x"40",
						   52598 => x"8A",		-- 00cd76: 8ACD            
						   52599 => x"CD",
						   -- Begin: __mspabi_srll
						   52600 => x"3E",		-- 00cd78: 3EF0             AND.W   #0x001f,R14
						   52601 => x"F0",
						   52602 => x"1F",		-- 00cd7a: 1F00            
						   52603 => x"00",
						   52604 => x"05",		-- 00cd7c: 0524             JEQ     (L_LSR_RET)
						   52605 => x"24",
						   -- Begin: L_LSR_TOP
						   52606 => x"12",		-- 00cd7e: 12C3             CLRC    
						   52607 => x"C3",
						   52608 => x"0D",		-- 00cd80: 0D10             RRC     R13
						   52609 => x"10",
						   52610 => x"0C",		-- 00cd82: 0C10             RRC     R12
						   52611 => x"10",
						   52612 => x"1E",		-- 00cd84: 1E83             DEC.W   R14
						   52613 => x"83",
						   52614 => x"FB",		-- 00cd86: FB23             JNE     (L_LSR_TOP)
						   52615 => x"23",
						   -- Begin: L_LSR_RET
						   52616 => x"30",		-- 00cd88: 3041             RET     
						   52617 => x"41",
						   -- Begin: memcpy
						   52618 => x"0E",		-- 00cd8a: 0E93             TST.W   R14
						   52619 => x"93",
						   52620 => x"06",		-- 00cd8c: 0624             JEQ     ($C$L2)
						   52621 => x"24",
						   52622 => x"0F",		-- 00cd8e: 0F4C             MOV.W   R12,R15
						   52623 => x"4C",
						   52624 => x"1F",		-- 00cd90: 1F53             INC.W   R15
						   52625 => x"53",
						   52626 => x"FF",		-- 00cd92: FF4D             MOV.B   @R13+,0xffff(R15)
						   52627 => x"4D",
						   52628 => x"FF",		-- 00cd94: FFFF            
						   52629 => x"FF",
						   52630 => x"1E",		-- 00cd96: 1E83             DEC.W   R14
						   52631 => x"83",
						   52632 => x"FB",		-- 00cd98: FB23             JNE     ($C$L1)
						   52633 => x"23",
						   52634 => x"30",		-- 00cd9a: 3041             RET     
						   52635 => x"41",
						   -- Begin: __mspabi_func_epilog_7
						   -- Begin: __mspabi_func_epilog
						   52636 => x"34",		-- 00cd9c: 3441             POP.W   R4
						   52637 => x"41",
						   -- Begin: __mspabi_func_epilog_6
						   52638 => x"35",		-- 00cd9e: 3541             POP.W   R5
						   52639 => x"41",
						   -- Begin: __mspabi_func_epilog_5
						   52640 => x"36",		-- 00cda0: 3641             POP.W   R6
						   52641 => x"41",
						   -- Begin: __mspabi_func_epilog_4
						   52642 => x"37",		-- 00cda2: 3741             POP.W   R7
						   52643 => x"41",
						   -- Begin: __mspabi_func_epilog_3
						   52644 => x"38",		-- 00cda4: 3841             POP.W   R8
						   52645 => x"41",
						   -- Begin: __mspabi_func_epilog_2
						   52646 => x"39",		-- 00cda6: 3941             POP.W   R9
						   52647 => x"41",
						   -- Begin: __mspabi_func_epilog_1
						   52648 => x"3A",		-- 00cda8: 3A41             POP.W   R10
						   52649 => x"41",
						   52650 => x"30",		-- 00cdaa: 3041             RET     
						   52651 => x"41",
						   -- Begin: strcpy
						   52652 => x"0F",		-- 00cdac: 0F4C             MOV.W   R12,R15
						   52653 => x"4C",
						   52654 => x"7E",		-- 00cdae: 7E4D             MOV.B   @R13+,R14
						   52655 => x"4D",
						   52656 => x"1F",		-- 00cdb0: 1F53             INC.W   R15
						   52657 => x"53",
						   52658 => x"CF",		-- 00cdb2: CF4E             MOV.B   R14,0xffff(R15)
						   52659 => x"4E",
						   52660 => x"FF",		-- 00cdb4: FFFF            
						   52661 => x"FF",
						   52662 => x"0E",		-- 00cdb6: 0E93             TST.W   R14
						   52663 => x"93",
						   52664 => x"FA",		-- 00cdb8: FA23             JNE     ($C$L1)
						   52665 => x"23",
						   52666 => x"30",		-- 00cdba: 3041             RET     
						   52667 => x"41",
						   -- Begin: strlen
						   52668 => x"3F",		-- 00cdbc: 3F43             MOV.W   #-1,R15
						   52669 => x"43",
						   52670 => x"1F",		-- 00cdbe: 1F53             INC.W   R15
						   52671 => x"53",
						   52672 => x"7E",		-- 00cdc0: 7E4C             MOV.B   @R12+,R14
						   52673 => x"4C",
						   52674 => x"0E",		-- 00cdc2: 0E93             TST.W   R14
						   52675 => x"93",
						   52676 => x"FC",		-- 00cdc4: FC23             JNE     ($C$L1)
						   52677 => x"23",
						   52678 => x"0C",		-- 00cdc6: 0C4F             MOV.W   R15,R12
						   52679 => x"4F",
						   52680 => x"30",		-- 00cdc8: 3041             RET     
						   52681 => x"41",
						   -- Begin: __mspabi_fltid
						   52682 => x"3C",		-- 00cdca: 3CB0             BIT.W   #0x8000,R12
						   52683 => x"B0",
						   52684 => x"00",		-- 00cdcc: 0080            
						   52685 => x"80",
						   52686 => x"0D",		-- 00cdce: 0D7D             SUBC.W  R13,R13
						   52687 => x"7D",
						   52688 => x"3D",		-- 00cdd0: 3DE3             INV.W   R13
						   52689 => x"E3",
						   52690 => x"30",		-- 00cdd2: 3040             BR      #__mspabi_fltlid
						   52691 => x"40",
						   52692 => x"B2",		-- 00cdd4: B2BA            
						   52693 => x"BA",
						   -- Begin: toupper
						   52694 => x"EC",		-- 00cdd6: ECB3             BIT.B   #2,0x8515(R12)
						   52695 => x"B3",
						   52696 => x"15",		-- 00cdd8: 1585            
						   52697 => x"85",
						   52698 => x"02",		-- 00cdda: 0224             JEQ     ($C$L1)
						   52699 => x"24",
						   52700 => x"3C",		-- 00cddc: 3C80             SUB.W   #0x0020,R12
						   52701 => x"80",
						   52702 => x"20",		-- 00cdde: 2000            
						   52703 => x"00",
						   52704 => x"30",		-- 00cde0: 3041             RET     
						   52705 => x"41",
						   -- Begin: abs
						   52706 => x"0C",		-- 00cde2: 0C93             TST.W   R12
						   52707 => x"93",
						   52708 => x"02",		-- 00cde4: 0234             JGE     ($C$L1)
						   52709 => x"34",
						   52710 => x"3C",		-- 00cde6: 3CE3             INV.W   R12
						   52711 => x"E3",
						   52712 => x"1C",		-- 00cde8: 1C53             INC.W   R12
						   52713 => x"53",
						   52714 => x"30",		-- 00cdea: 3041             RET     
						   52715 => x"41",
						   -- Begin: malloc
						   52716 => x"0D",		-- 00cdec: 0D4C             MOV.W   R12,R13
						   52717 => x"4C",
						   52718 => x"2C",		-- 00cdee: 2C42             MOV.W   #4,R12
						   52719 => x"42",
						   52720 => x"30",		-- 00cdf0: 3040             BR      #aligned_alloc
						   52721 => x"40",
						   52722 => x"00",		-- 00cdf2: 00B4            
						   52723 => x"B4",
						   -- Begin: _outc
						   52724 => x"4C",		-- 00cdf4: 4C4C             MOV.B   R12,R12
						   52725 => x"4C",
						   52726 => x"30",		-- 00cdf6: 3040             BR      #fputc
						   52727 => x"40",
						   52728 => x"9C",		-- 00cdf8: 9CBC            
						   52729 => x"BC",
						   -- Begin: abort
						   52730 => x"03",		-- 00cdfa: 0343             NOP     
						   52731 => x"43",
						   52732 => x"FF",		-- 00cdfc: FF3F             JMP     ($C$L1)
						   52733 => x"3F",
						   52734 => x"03",		-- 00cdfe: 0343             NOP     
						   52735 => x"43",
						   -- Begin: _outs
						   52736 => x"30",		-- 00ce00: 3040             BR      #fputs
						   52737 => x"40",
						   52738 => x"F6",		-- 00ce02: F6B4            
						   52739 => x"B4",
						   -- Begin: _system_pre_init
						   52740 => x"1C",		-- 00ce04: 1C43             MOV.W   #1,R12
						   52741 => x"43",
						   52742 => x"30",		-- 00ce06: 3041             RET     
						   52743 => x"41",
						   -- Begin: _nop
						   52744 => x"30",		-- 00ce08: 3041             RET     
						   52745 => x"41",
						   -- Begin: _system_post_cinit
						   52746 => x"30",		-- 00ce0a: 3041             RET     
						   52747 => x"41",
						   -- ISR Trap
						   52748 => x"32",		-- 00ce0c: 32D0             BIS.W   #0x0010,SR
						   52749 => x"D0",
						   52750 => x"10",		-- 00ce0e: 1000            
						   52751 => x"00",
						   52752 => x"FD",		-- 00ce10: FD3F             JMP     (__TI_ISR_TRAP)
						   52753 => x"3F",
						   52754 => x"03",		-- 00ce12: 0343             NOP     
						   52755 => x"43",
						   -- IRQ Vectors (Interrupt Vectors)
						   65486 => x"0c",		-- 00ffce:ce0c PORT4 __TI_int22 int22
						   65487 => x"ce",
						   65488 => x"0c",		-- 00ffd0:ce0c PORT3 __TI_int23 int23
						   65489 => x"ce",
						   65490 => x"0c",		-- 00ffd2:ce0c PORT2 __TI_int24 int24
						   65491 => x"ce",
						   65492 => x"0c",		-- 00ffd4:ce0c PORT1 __TI_int25 int25
						   65493 => x"ce",
						   65494 => x"0c",		-- 00ffd6:ce0c SAC1_SAC3 __TI_int26 int26
						   65495 => x"ce",
						   65496 => x"0c",		-- 00ffd8:ce0c SAC0_SAC2 __TI_int27 int27
						   65497 => x"ce",
						   65498 => x"0c",		-- 00ffda:ce0c ECOMP0_ECOMP1 __TI_int28 int28
						   65499 => x"ce",
						   65500 => x"0c",		-- 00ffdc:ce0c ADC __TI_int29 int29
						   65501 => x"ce",
						   65502 => x"0c",		-- 00ffde:ce0c EUSCI_B1 __TI_int30 int30
						   65503 => x"ce",
						   65504 => x"0c",		-- 00ffe0:ce0c EUSCI_B0 __TI_int31 int31
						   65505 => x"ce",
						   65506 => x"0c",		-- 00ffe2:ce0c EUSCI_A1 __TI_int32 int32
						   65507 => x"ce",
						   65508 => x"0c",		-- 00ffe4:ce0c EUSCI_A0 __TI_int33 int33
						   65509 => x"ce",
						   65510 => x"0c",		-- 00ffe6:ce0c WDT __TI_int34 int34
						   65511 => x"ce",
						   65512 => x"0c",		-- 00ffe8:ce0c RTC __TI_int35 int35
						   65513 => x"ce",
						   65514 => x"0c",		-- 00ffea:ce0c TIMER3_B1 __TI_int36 int36
						   65515 => x"ce",
						   65516 => x"0c",		-- 00ffec:ce0c TIMER3_B0 __TI_int37 int37
						   65517 => x"ce",
						   65518 => x"0c",		-- 00ffee:ce0c TIMER2_B1 __TI_int38 int38
						   65519 => x"ce",
						   65520 => x"0c",		-- 00fff0:ce0c TIMER2_B0 __TI_int39 int39
						   65521 => x"ce",
						   65522 => x"0c",		-- 00fff2:ce0c TIMER1_B1 __TI_int40 int40
						   65523 => x"ce",
						   65524 => x"0c",		-- 00fff4:ce0c TIMER1_B0 __TI_int41 int41
						   65525 => x"ce",
						   65526 => x"0c",		-- 00fff6:ce0c TIMER0_B1 __TI_int42 int42
						   65527 => x"ce",
						   65528 => x"0c",		-- 00fff8:ce0c TIMER0_B0 __TI_int43 int43
						   65529 => x"ce",
						   65530 => x"0c",		-- 00fffa:ce0c UNMI __TI_int44 int44
						   65531 => x"ce",
						   65532 => x"0c",		-- 00fffc:ce0c SYSNMI __TI_int45 int45
						   65533 => x"ce",

                           65534 =>  x"00",		-- Reset Vector = xFFFE:xFFFF
                           65535 =>  x"80",		--  Startup Value = x8000

                           others => x"00");

    signal EN : std_logic;
    
    begin
    -- Note 1:  The bus system uses a 16-bit Address (MAB)
    --          This address size can access locations from x0000 to xFFFF
    --          But our array is only defined from x8000 to xFFFF and
    --          if we try to access it with any other address, it will crash.
    --          So the first thing we need to do is create a local enable that
    --          will only assert when MAB is within x8000 to xFFFF.

     LOCAL_EN : process (MAB) 
     begin
         if ( (to_integer(unsigned(MAB)) >= 32768) and (to_integer(unsigned(MAB)) <= 65535)) then
           EN <= '1';
         else 
           EN <= '0';
         end if;
     end process;

    
    -- Note 2:  The bus system uses a 16-bit Address (MAB)
    --          The MDB_out is also provided as a 16-bit word
    --          However, the memory array is actually built as 8-bit bytes.
    --          So for a given 16-bit MAB, we give MDB_out = HB : LB
    --                                                 or  = ROM(MAB);1) : ROM(MAB)

    MEMORY_ROM : process (clk) 
    begin
        if (rising_edge(clk)) then
            if (EN='1' and write='0') then                      
              MDB_in <= ROM(to_integer(unsigned(MAB)) + 1 ) & ROM(to_integer(unsigned(MAB))); 
            end if;
        end if;
    end process;


end architecture;