library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;


entity highroller_memory is
    port ( clk	: in	std_logic;
         MAB		: in	std_logic_vector(15 downto 0);
         MDB_in  	: out	std_logic_vector(15 downto 0);
         MDB_out  	: in	std_logic_vector(15 downto 0);
         write	    : in	std_logic;
         Byte       : in    std_logic);
end entity;

architecture highroller_memory_arch of highroller_memory is

type rom_type is array (32768 to 65535) of std_logic_vector(7 downto 0);  -- this is MAB: x8000 to xFFFF
    
constant ROM : rom_type :=(32768 => x"00",		-- Begin: .cinit DATA Section
						   32769 => x"ff",
						   32770 => x"00",
						   32771 => x"38",
						   32772 => x"28",
						   32773 => x"37",
						   32774 => x"18",
						   32775 => x"00",
						   32776 => x"27",
						   32777 => x"34",
						   32778 => x"ff",
						   32779 => x"08",
						   32780 => x"39",
						   32781 => x"00",
						   32782 => x"00",
						   32783 => x"17",
						   32784 => x"00",
						   32785 => x"24",
						   32786 => x"0d",
						   32787 => x"ff",
						   32788 => x"78",
						   32789 => x"00",
						   32790 => x"29",
						   32791 => x"36",
						   32794 => x"00",
						   32795 => x"35",
						   32796 => x"fd",
						   32797 => x"07",
						   32798 => x"00",
						   32799 => x"40",
						   32800 => x"14",
						   32801 => x"13",
						   32802 => x"7d",
						   32803 => x"12",
						   32804 => x"68",
						   32805 => x"69",
						   32806 => x"ff",
						   32807 => x"00",
						   32808 => x"00",
						   32809 => x"19",
						   32810 => x"6a",
						   32811 => x"26",
						   32814 => x"3a",
						   32815 => x"be",
						   32816 => x"01",
						   32817 => x"50",
						   32818 => x"00",
						   32819 => x"25",
						   32820 => x"0e",
						   32821 => x"77",
						   32822 => x"76",
						   32823 => x"01",
						   32824 => x"d0",
						   32825 => x"6b",
						   32826 => x"ff",
						   32827 => x"00",
						   32828 => x"00",
						   32829 => x"04",
						   32830 => x"00",
						   32831 => x"03",
						   32832 => x"00",
						   32833 => x"6d",
						   32834 => x"6c",
						   32835 => x"df",
						   32836 => x"02",
						   32837 => x"01",
						   32838 => x"58",
						   32839 => x"00",
						   32840 => x"59",
						   32841 => x"01",
						   32842 => x"81",
						   32843 => x"33",
						   32844 => x"09",
						   32845 => x"ff",
						   32846 => x"0a",
						   32847 => x"5a",
						   32848 => x"00",
						   32849 => x"16",
						   32850 => x"0b",
						   32851 => x"00",
						   32852 => x"0c",
						   32853 => x"00",
						   32854 => x"e7",
						   32855 => x"00",
						   32856 => x"2a",
						   32857 => x"2b",
						   32858 => x"02",
						   32859 => x"91",
						   32860 => x"02",
						   32861 => x"d1",
						   32862 => x"15",
						   32863 => x"00",
						   32864 => x"7e",
						   32865 => x"af",
						   32866 => x"7f",
						   32867 => x"67",
						   32868 => x"00",
						   32869 => x"66",
						   32870 => x"00",
						   32871 => x"e4",
						   32872 => x"5b",
						   32873 => x"01",
						   32874 => x"62",
						   32875 => x"74",
						   32876 => x"ef",
						   32877 => x"75",
						   32880 => x"73",
						   32881 => x"06",
						   32882 => x"00",
						   32883 => x"5d",
						   32884 => x"5e",
						   32885 => x"5c",
						   32886 => x"ff",
						   32887 => x"00",
						   32888 => x"72",
						   32889 => x"5f",
						   32890 => x"71",
						   32891 => x"00",
						   32892 => x"48",
						   32893 => x"47",
						   32894 => x"00",
						   32895 => x"ff",
						   32896 => x"44",
						   32897 => x"49",
						   32900 => x"1d",
						   32901 => x"00",
						   32902 => x"46",
						   32903 => x"00",
						   32904 => x"ff",
						   32905 => x"45",
						   32908 => x"23",
						   32909 => x"22",
						   32910 => x"79",
						   32911 => x"00",
						   32912 => x"7a",
						   32913 => x"ff",
						   32914 => x"00",
						   32915 => x"4a",
						   32918 => x"1e",
						   32919 => x"06",
						   32920 => x"00",
						   32921 => x"7b",
						   32922 => x"f6",
						   32923 => x"08",
						   32924 => x"60",
						   32925 => x"7c",
						   32926 => x"11",
						   32927 => x"08",
						   32928 => x"b0",
						   32929 => x"43",
						   32930 => x"1a",
						   32931 => x"00",
						   32932 => x"1b",
						   32933 => x"57",
						   32934 => x"1c",
						   32935 => x"00",
						   32936 => x"3b",
						   32937 => x"05",
						   32938 => x"52",
						   32939 => x"0f",
						   32940 => x"05",
						   32941 => x"b5",
						   32942 => x"05",
						   32943 => x"0a",
						   32944 => x"40",
						   32945 => x"ff",
						   32946 => x"6e",
						   32947 => x"00",
						   32948 => x"6f",
						   32949 => x"10",
						   32950 => x"57",
						   32951 => x"54",
						   32952 => x"00",
						   32953 => x"2d",
						   32954 => x"af",
						   32955 => x"56",
						   32956 => x"55",
						   32957 => x"00",
						   32958 => x"32",
						   32959 => x"0b",
						   32960 => x"30",
						   32961 => x"2e",
						   32962 => x"0b",
						   32963 => x"70",
						   32964 => x"21",
						   32965 => x"ff",
						   32966 => x"00",
						   32967 => x"53",
						   32968 => x"00",
						   32969 => x"2c",
						   32970 => x"4b",
						   32971 => x"00",
						   32972 => x"00",
						   32973 => x"1f",
						   32974 => x"fe",
						   32975 => x"08",
						   32976 => x"34",
						   32977 => x"20",
						   32978 => x"64",
						   32979 => x"3d",
						   32980 => x"65",
						   32981 => x"42",
						   32982 => x"00",
						   32983 => x"3e",
						   32984 => x"bf",
						   32985 => x"00",
						   32986 => x"31",
						   32987 => x"63",
						   32988 => x"3c",
						   32989 => x"00",
						   32990 => x"2f",
						   32991 => x"0d",
						   32992 => x"70",
						   32993 => x"30",
						   32994 => x"ff",
						   32995 => x"4d",
						   32996 => x"52",
						   32997 => x"4e",
						   32998 => x"41",
						   32999 => x"4c",
						   33000 => x"3f",
						   33001 => x"00",
						   33002 => x"40",
						   33003 => x"ff",
						   33004 => x"62",
						   33005 => x"51",
						   33006 => x"4f",
						   33007 => x"50",
						   33008 => x"61",
						   33009 => x"60",
						   33010 => x"70",
						   33011 => x"00",
						   33012 => x"0f",
						   33013 => x"e8",
						   33014 => x"03",
						   33015 => x"3d",
						   33016 => x"00",
						   33017 => x"ff",
						   33018 => x"f0",
						   33019 => x"00",
						   33020 => x"c6",
						   33021 => x"81",
						   33022 => x"2a",
						   33023 => x"83",
						   33024 => x"00",
						   33025 => x"80",
						   33026 => x"00",
						   33027 => x"20",
						   -- Begin: program memory TEXT Section
						   33028 => x"21",		-- 008104: 2183             DECD.W  SP
						   33029 => x"A3",
						   33030 => x"B2",		-- 008106: B240             MOV.W   #0x5a80,&WDTCTL_L
						   33031 => x"60",
						   33032 => x"80",		-- 008108: 805A            
						   33033 => x"5A",
						   33034 => x"CC",		-- 00810a: CC01            
						   33035 => x"01",
						   33036 => x"92",		-- 00810c: 92C3             BIC.W   #1,&PM5CTL0_L
						   33037 => x"E3",
						   33038 => x"30",		-- 00810e: 3001            
						   33039 => x"01",
						   33040 => x"5F",		-- 008110: 5F42             MOV.B   &P1DIR,R15
						   33041 => x"62",
						   33042 => x"04",		-- 008112: 0402            
						   33043 => x"02",
						   33044 => x"C2",		-- 008114: C243             CLR.B   &P1DIR
						   33045 => x"63",
						   33046 => x"04",		-- 008116: 0402            
						   33047 => x"02",
						   33048 => x"F2",		-- 008118: F2F0             AND.B   #0x00fc,&P2DIR
						   33049 => x"10",
						   33050 => x"FC",		-- 00811a: FC00            
						   33051 => x"00",
						   33052 => x"05",		-- 00811c: 0502            
						   33053 => x"02",
						   33054 => x"F2",		-- 00811e: F2D0             BIS.B   #0x0034,&P2DIR
						   33055 => x"F0",
						   33056 => x"34",		-- 008120: 3400            
						   33057 => x"00",
						   33058 => x"05",		-- 008122: 0502            
						   33059 => x"02",
						   33060 => x"B2",		-- 008124: B2D0             BIS.W   #0x0220,&TB0CTL_L
						   33061 => x"F0",
						   33062 => x"20",		-- 008126: 2002            
						   33063 => x"02",
						   33064 => x"80",		-- 008128: 8003            
						   33065 => x"03",
						   33066 => x"B2",		-- 00812a: B2D0             BIS.W   #0x0010,&TB0CCTL0_L
						   33067 => x"F0",
						   33068 => x"10",		-- 00812c: 1000            
						   33069 => x"00",
						   33070 => x"82",		-- 00812e: 8203            
						   33071 => x"03",
						   33072 => x"92",		-- 008130: 9242             MOV.W   &frequency,&TB0CCR0_L
						   33073 => x"62",
						   33074 => x"00",		-- 008132: 0021            
						   33075 => x"21",
						   33076 => x"92",		-- 008134: 9203            
						   33077 => x"03",
						   33078 => x"32",		-- 008136: 32D2             EINT    
						   33079 => x"F2",
						   33080 => x"92",		-- 008138: 92D3             BIS.W   #1,&UCA1IE_L
						   33081 => x"F3",
						   33082 => x"9A",		-- 00813a: 9A05            
						   33083 => x"05",
						   33084 => x"3F",		-- 00813c: 3F40             MOV.W   #0x0003,R15
						   33085 => x"60",
						   33086 => x"03",		-- 00813e: 0300            
						   33087 => x"00",
						   33088 => x"5F",		-- 008140: 5FF2             AND.B   &P2IN,R15
						   33089 => x"12",
						   33090 => x"01",		-- 008142: 0102            
						   33091 => x"02",
						   33092 => x"C1",		-- 008144: C14F             MOV.B   R15,0x0000(SP)
						   33093 => x"6F",
						   33094 => x"00",		-- 008146: 0000            
						   33095 => x"00",
						   33096 => x"D1",		-- 008148: D193             CMP.B   #1,0x0000(SP)
						   33097 => x"B3",
						   33098 => x"00",		-- 00814a: 0000            
						   33099 => x"00",
						   33100 => x"04",		-- 00814c: 0420             JNE     ($C$L2)
						   33101 => x"40",
						   33102 => x"B2",		-- 00814e: B240             MOV.W   #0x002f,&set_angle
						   33103 => x"60",
						   33104 => x"2F",		-- 008150: 2F00            
						   33105 => x"00",
						   33106 => x"02",		-- 008152: 0221            
						   33107 => x"21",
						   33108 => x"0A",		-- 008154: 0A3C             JMP     ($C$L4)
						   33109 => x"5C",
						   33110 => x"E1",		-- 008156: E193             CMP.B   #2,0x0000(SP)
						   33111 => x"B3",
						   33112 => x"00",		-- 008158: 0000            
						   33113 => x"00",
						   33114 => x"04",		-- 00815a: 0420             JNE     ($C$L3)
						   33115 => x"40",
						   33116 => x"B2",		-- 00815c: B240             MOV.W   #0x004f,&set_angle
						   33117 => x"60",
						   33118 => x"4F",		-- 00815e: 4F00            
						   33119 => x"00",
						   33120 => x"02",		-- 008160: 0221            
						   33121 => x"21",
						   33122 => x"03",		-- 008162: 033C             JMP     ($C$L4)
						   33123 => x"5C",
						   33124 => x"B2",		-- 008164: B240             MOV.W   #0x003d,&set_angle
						   33125 => x"60",
						   33126 => x"3D",		-- 008166: 3D00            
						   33127 => x"00",
						   33128 => x"02",		-- 008168: 0221            
						   33129 => x"21",
						   33130 => x"5F",		-- 00816a: 5F42             MOV.B   &P1IN,R15
						   33131 => x"62",
						   33132 => x"00",		-- 00816c: 0002            
						   33133 => x"02",
						   33134 => x"D1",		-- 00816e: D14F             MOV.B   0x2000(R15),0x0000(SP)
						   33135 => x"6F",
						   33136 => x"00",		-- 008170: 0020            
						   33137 => x"20",
						   33138 => x"00",		-- 008172: 0000            
						   33139 => x"00",
						   33140 => x"6F",		-- 008174: 6F41             MOV.B   @SP,R15
						   33141 => x"61",
						   33142 => x"1F",		-- 008176: 1F92             CMP.W   &set_angle,R15
						   33143 => x"B2",
						   33144 => x"02",		-- 008178: 0221            
						   33145 => x"21",
						   33146 => x"0B",		-- 00817a: 0B2C             JHS     ($C$L5)
						   33147 => x"4C",
						   33148 => x"E2",		-- 00817c: E2C2             BIC.B   #4,&P2OUT
						   33149 => x"E2",
						   33150 => x"03",		-- 00817e: 0302            
						   33151 => x"02",
						   33152 => x"F2",		-- 008180: F2F0             AND.B   #0x00df,&P2OUT
						   33153 => x"10",
						   33154 => x"DF",		-- 008182: DF00            
						   33155 => x"00",
						   33156 => x"03",		-- 008184: 0302            
						   33157 => x"02",
						   33158 => x"5F",		-- 008186: 5F42             MOV.B   &set_angle,R15
						   33159 => x"62",
						   33160 => x"02",		-- 008188: 0221            
						   33161 => x"21",
						   33162 => x"6F",		-- 00818a: 6F81             SUB.B   @SP,R15
						   33163 => x"A1",
						   33164 => x"C1",		-- 00818c: C14F             MOV.B   R15,0x0000(SP)
						   33165 => x"6F",
						   33166 => x"00",		-- 00818e: 0000            
						   33167 => x"00",
						   33168 => x"0F",		-- 008190: 0F3C             JMP     ($C$L7)
						   33169 => x"5C",
						   33170 => x"6F",		-- 008192: 6F41             MOV.B   @SP,R15
						   33171 => x"61",
						   33172 => x"82",		-- 008194: 829F             CMP.W   R15,&set_angle
						   33173 => x"BF",
						   33174 => x"02",		-- 008196: 0221            
						   33175 => x"21",
						   33176 => x"09",		-- 008198: 092C             JHS     ($C$L6)
						   33177 => x"4C",
						   33178 => x"E2",		-- 00819a: E2C2             BIC.B   #4,&P2OUT
						   33179 => x"E2",
						   33180 => x"03",		-- 00819c: 0302            
						   33181 => x"02",
						   33182 => x"F2",		-- 00819e: F2D0             BIS.B   #0x0020,&P2OUT
						   33183 => x"F0",
						   33184 => x"20",		-- 0081a0: 2000            
						   33185 => x"00",
						   33186 => x"03",		-- 0081a2: 0302            
						   33187 => x"02",
						   33188 => x"D1",		-- 0081a4: D182             SUB.B   &set_angle,0x0000(SP)
						   33189 => x"A2",
						   33190 => x"02",		-- 0081a6: 0221            
						   33191 => x"21",
						   33192 => x"00",		-- 0081a8: 0000            
						   33193 => x"00",
						   33194 => x"02",		-- 0081aa: 023C             JMP     ($C$L7)
						   33195 => x"5C",
						   33196 => x"E2",		-- 0081ac: E2D2             BIS.B   #4,&P2OUT
						   33197 => x"F2",
						   33198 => x"03",		-- 0081ae: 0302            
						   33199 => x"02",
						   33200 => x"6F",		-- 0081b0: 6F41             MOV.B   @SP,R15
						   33201 => x"61",
						   33202 => x"0C",		-- 0081b2: 0C4F             MOV.W   R15,R12
						   33203 => x"6F",
						   33204 => x"B0",		-- 0081b4: B012             CALL    #__mspabi_slli_6
						   33205 => x"32",
						   33206 => x"EE",		-- 0081b6: EE82            
						   33207 => x"82",
						   33208 => x"0C",		-- 0081b8: 0C8F             SUB.W   R15,R12
						   33209 => x"AF",
						   33210 => x"3F",		-- 0081ba: 3F40             MOV.W   #0x0fa0,R15
						   33211 => x"60",
						   33212 => x"A0",		-- 0081bc: A00F            
						   33213 => x"0F",
						   33214 => x"0F",		-- 0081be: 0F8C             SUB.W   R12,R15
						   33215 => x"AC",
						   33216 => x"82",		-- 0081c0: 824F             MOV.W   R15,&frequency
						   33217 => x"6F",
						   33218 => x"00",		-- 0081c2: 0021            
						   33219 => x"21",
						   33220 => x"BB",		-- 0081c4: BB3F             JMP     ($C$L1)
						   33221 => x"5F",
						   -- Begin: __TI_decompress_lzss
						   33222 => x"0A",		-- 0081c6: 0A12             PUSH    R10
						   33223 => x"32",
						   33224 => x"09",		-- 0081c8: 0912             PUSH    R9
						   33225 => x"32",
						   33226 => x"08",		-- 0081ca: 0812             PUSH    R8
						   33227 => x"32",
						   33228 => x"0A",		-- 0081cc: 0A4C             MOV.W   R12,R10
						   33229 => x"6C",
						   33230 => x"78",		-- 0081ce: 784A             MOV.B   @R10+,R8
						   33231 => x"6A",
						   33232 => x"09",		-- 0081d0: 0943             CLR.W   R9
						   33233 => x"63",
						   33234 => x"11",		-- 0081d2: 113C             JMP     ($C$L6)
						   33235 => x"5C",
						   33236 => x"0E",		-- 0081d4: 0E4D             MOV.W   R13,R14
						   33237 => x"6D",
						   33238 => x"0E",		-- 0081d6: 0E8B             SUB.W   R11,R14
						   33239 => x"AB",
						   33240 => x"1E",		-- 0081d8: 1E83             DEC.W   R14
						   33241 => x"A3",
						   33242 => x"1D",		-- 0081da: 1D53             INC.W   R13
						   33243 => x"73",
						   33244 => x"FD",		-- 0081dc: FD4E             MOV.B   @R14+,0xffff(R13)
						   33245 => x"6E",
						   33246 => x"FF",		-- 0081de: FFFF            
						   33247 => x"FF",
						   33248 => x"1F",		-- 0081e0: 1F83             DEC.W   R15
						   33249 => x"A3",
						   33250 => x"FB",		-- 0081e2: FB23             JNE     ($C$L3)
						   33251 => x"43",
						   33252 => x"03",		-- 0081e4: 033C             JMP     ($C$L5)
						   33253 => x"5C",
						   33254 => x"1D",		-- 0081e6: 1D53             INC.W   R13
						   33255 => x"73",
						   33256 => x"FD",		-- 0081e8: FD4A             MOV.B   @R10+,0xffff(R13)
						   33257 => x"6A",
						   33258 => x"FF",		-- 0081ea: FFFF            
						   33259 => x"FF",
						   33260 => x"12",		-- 0081ec: 12C3             CLRC    
						   33261 => x"E3",
						   33262 => x"08",		-- 0081ee: 0810             RRC     R8
						   33263 => x"30",
						   33264 => x"19",		-- 0081f0: 1953             INC.W   R9
						   33265 => x"73",
						   33266 => x"39",		-- 0081f2: 3992             CMP.W   #8,R9
						   33267 => x"B2",
						   33268 => x"EC",		-- 0081f4: EC37             JGE     ($C$L1)
						   33269 => x"57",
						   33270 => x"18",		-- 0081f6: 18B3             BIT.W   #1,R8
						   33271 => x"D3",
						   33272 => x"F6",		-- 0081f8: F623             JNE     ($C$L4)
						   33273 => x"43",
						   33274 => x"7B",		-- 0081fa: 7B4A             MOV.B   @R10+,R11
						   33275 => x"6A",
						   33276 => x"7F",		-- 0081fc: 7F4A             MOV.B   @R10+,R15
						   33277 => x"6A",
						   33278 => x"0C",		-- 0081fe: 0C4B             MOV.W   R11,R12
						   33279 => x"6B",
						   33280 => x"B0",		-- 008200: B012             CALL    #__mspabi_slli_4
						   33281 => x"32",
						   33282 => x"F2",		-- 008202: F282            
						   33283 => x"82",
						   33284 => x"0B",		-- 008204: 0B4C             MOV.W   R12,R11
						   33285 => x"6C",
						   33286 => x"0C",		-- 008206: 0C4F             MOV.W   R15,R12
						   33287 => x"6F",
						   33288 => x"B0",		-- 008208: B012             CALL    #__mspabi_srli_4
						   33289 => x"32",
						   33290 => x"7C",		-- 00820a: 7C82            
						   33291 => x"82",
						   33292 => x"3C",		-- 00820c: 3CF0             AND.W   #0x000f,R12
						   33293 => x"10",
						   33294 => x"0F",		-- 00820e: 0F00            
						   33295 => x"00",
						   33296 => x"0B",		-- 008210: 0BDC             BIS.W   R12,R11
						   33297 => x"FC",
						   33298 => x"3F",		-- 008212: 3FF0             AND.W   #0x000f,R15
						   33299 => x"10",
						   33300 => x"0F",		-- 008214: 0F00            
						   33301 => x"00",
						   33302 => x"3F",		-- 008216: 3F50             ADD.W   #0x0003,R15
						   33303 => x"70",
						   33304 => x"03",		-- 008218: 0300            
						   33305 => x"00",
						   33306 => x"3F",		-- 00821a: 3F90             CMP.W   #0x0012,R15
						   33307 => x"B0",
						   33308 => x"12",		-- 00821c: 1200            
						   33309 => x"00",
						   33310 => x"0C",		-- 00821e: 0C20             JNE     ($C$L8)
						   33311 => x"40",
						   33312 => x"7E",		-- 008220: 7E4A             MOV.B   @R10+,R14
						   33313 => x"6A",
						   33314 => x"3E",		-- 008222: 3EB0             BIT.W   #0x0080,R14
						   33315 => x"D0",
						   33316 => x"80",		-- 008224: 8000            
						   33317 => x"00",
						   33318 => x"07",		-- 008226: 0724             JEQ     ($C$L7)
						   33319 => x"44",
						   33320 => x"7C",		-- 008228: 7C4A             MOV.B   @R10+,R12
						   33321 => x"6A",
						   33322 => x"4C",		-- 00822a: 4C4C             MOV.B   R12,R12
						   33323 => x"6C",
						   33324 => x"B0",		-- 00822c: B012             CALL    #__mspabi_slli_7
						   33325 => x"32",
						   33326 => x"EC",		-- 00822e: EC82            
						   33327 => x"82",
						   33328 => x"3E",		-- 008230: 3EF0             AND.W   #0x007f,R14
						   33329 => x"10",
						   33330 => x"7F",		-- 008232: 7F00            
						   33331 => x"00",
						   33332 => x"0E",		-- 008234: 0EDC             BIS.W   R12,R14
						   33333 => x"FC",
						   33334 => x"0F",		-- 008236: 0F5E             ADD.W   R14,R15
						   33335 => x"7E",
						   33336 => x"3B",		-- 008238: 3B90             CMP.W   #0x0fff,R11
						   33337 => x"B0",
						   33338 => x"FF",		-- 00823a: FF0F            
						   33339 => x"0F",
						   33340 => x"CB",		-- 00823c: CB23             JNE     ($C$L2)
						   33341 => x"43",
						   33342 => x"30",		-- 00823e: 3040             BR      #__mspabi_func_epilog_3
						   33343 => x"60",
						   33344 => x"56",		-- 008240: 5683            
						   33345 => x"83",
						   -- Begin: __mspabi_srli
						   33346 => x"3D",		-- 008242: 3DF0             AND.W   #0x000f,R13
						   33347 => x"10",
						   33348 => x"0F",		-- 008244: 0F00            
						   33349 => x"00",
						   33350 => x"3D",		-- 008246: 3DE0             XOR.W   #0x000f,R13
						   33351 => x"00",
						   33352 => x"0F",		-- 008248: 0F00            
						   33353 => x"00",
						   33354 => x"0D",		-- 00824a: 0D5D             RLA.W   R13
						   33355 => x"7D",
						   33356 => x"0D",		-- 00824c: 0D5D             RLA.W   R13
						   33357 => x"7D",
						   33358 => x"00",		-- 00824e: 005D             ADD.W   R13,PC
						   33359 => x"7D",
						   -- Begin: __mspabi_srli_15
						   33360 => x"12",		-- 008250: 12C3             CLRC    
						   33361 => x"E3",
						   33362 => x"0C",		-- 008252: 0C10             RRC     R12
						   33363 => x"30",
						   -- Begin: __mspabi_srli_14
						   33364 => x"12",		-- 008254: 12C3             CLRC    
						   33365 => x"E3",
						   33366 => x"0C",		-- 008256: 0C10             RRC     R12
						   33367 => x"30",
						   -- Begin: __mspabi_srli_13
						   33368 => x"12",		-- 008258: 12C3             CLRC    
						   33369 => x"E3",
						   33370 => x"0C",		-- 00825a: 0C10             RRC     R12
						   33371 => x"30",
						   -- Begin: __mspabi_srli_12
						   33372 => x"12",		-- 00825c: 12C3             CLRC    
						   33373 => x"E3",
						   33374 => x"0C",		-- 00825e: 0C10             RRC     R12
						   33375 => x"30",
						   -- Begin: __mspabi_srli_11
						   33376 => x"12",		-- 008260: 12C3             CLRC    
						   33377 => x"E3",
						   33378 => x"0C",		-- 008262: 0C10             RRC     R12
						   33379 => x"30",
						   -- Begin: __mspabi_srli_10
						   33380 => x"12",		-- 008264: 12C3             CLRC    
						   33381 => x"E3",
						   33382 => x"0C",		-- 008266: 0C10             RRC     R12
						   33383 => x"30",
						   -- Begin: __mspabi_srli_9
						   33384 => x"12",		-- 008268: 12C3             CLRC    
						   33385 => x"E3",
						   33386 => x"0C",		-- 00826a: 0C10             RRC     R12
						   33387 => x"30",
						   -- Begin: __mspabi_srli_8
						   33388 => x"12",		-- 00826c: 12C3             CLRC    
						   33389 => x"E3",
						   33390 => x"0C",		-- 00826e: 0C10             RRC     R12
						   33391 => x"30",
						   -- Begin: __mspabi_srli_7
						   33392 => x"12",		-- 008270: 12C3             CLRC    
						   33393 => x"E3",
						   33394 => x"0C",		-- 008272: 0C10             RRC     R12
						   33395 => x"30",
						   -- Begin: __mspabi_srli_6
						   33396 => x"12",		-- 008274: 12C3             CLRC    
						   33397 => x"E3",
						   33398 => x"0C",		-- 008276: 0C10             RRC     R12
						   33399 => x"30",
						   -- Begin: __mspabi_srli_5
						   33400 => x"12",		-- 008278: 12C3             CLRC    
						   33401 => x"E3",
						   33402 => x"0C",		-- 00827a: 0C10             RRC     R12
						   33403 => x"30",
						   -- Begin: __mspabi_srli_4
						   33404 => x"12",		-- 00827c: 12C3             CLRC    
						   33405 => x"E3",
						   33406 => x"0C",		-- 00827e: 0C10             RRC     R12
						   33407 => x"30",
						   -- Begin: __mspabi_srli_3
						   33408 => x"12",		-- 008280: 12C3             CLRC    
						   33409 => x"E3",
						   33410 => x"0C",		-- 008282: 0C10             RRC     R12
						   33411 => x"30",
						   -- Begin: __mspabi_srli_2
						   33412 => x"12",		-- 008284: 12C3             CLRC    
						   33413 => x"E3",
						   33414 => x"0C",		-- 008286: 0C10             RRC     R12
						   33415 => x"30",
						   -- Begin: __mspabi_srli_1
						   33416 => x"12",		-- 008288: 12C3             CLRC    
						   33417 => x"E3",
						   33418 => x"0C",		-- 00828a: 0C10             RRC     R12
						   33419 => x"30",
						   33420 => x"30",		-- 00828c: 3041             RET     
						   33421 => x"61",
						   -- Begin: __TI_auto_init_nobinit_nopinit
						   33422 => x"0A",		-- 00828e: 0A12             PUSH    R10
						   33423 => x"32",
						   33424 => x"09",		-- 008290: 0912             PUSH    R9
						   33425 => x"32",
						   33426 => x"3F",		-- 008292: 3F40             MOV.W   #0x80fc,R15
						   33427 => x"60",
						   33428 => x"FC",		-- 008294: FC80            
						   33429 => x"80",
						   33430 => x"3F",		-- 008296: 3F90             CMP.W   #0x8100,R15
						   33431 => x"B0",
						   33432 => x"00",		-- 008298: 0081            
						   33433 => x"81",
						   33434 => x"16",		-- 00829a: 1624             JEQ     ($C$L22)
						   33435 => x"44",
						   33436 => x"3F",		-- 00829c: 3F40             MOV.W   #0x8100,R15
						   33437 => x"60",
						   33438 => x"00",		-- 00829e: 0081            
						   33439 => x"81",
						   33440 => x"3F",		-- 0082a0: 3F90             CMP.W   #0x8104,R15
						   33441 => x"B0",
						   33442 => x"04",		-- 0082a2: 0481            
						   33443 => x"81",
						   33444 => x"11",		-- 0082a4: 1124             JEQ     ($C$L22)
						   33445 => x"44",
						   33446 => x"3A",		-- 0082a6: 3A40             MOV.W   #0x8104,R10
						   33447 => x"60",
						   33448 => x"04",		-- 0082a8: 0481            
						   33449 => x"81",
						   33450 => x"3A",		-- 0082aa: 3A80             SUB.W   #0x8100,R10
						   33451 => x"A0",
						   33452 => x"00",		-- 0082ac: 0081            
						   33453 => x"81",
						   33454 => x"0A",		-- 0082ae: 0A11             RRA     R10
						   33455 => x"31",
						   33456 => x"0A",		-- 0082b0: 0A11             RRA     R10
						   33457 => x"31",
						   33458 => x"39",		-- 0082b2: 3940             MOV.W   #0x8100,R9
						   33459 => x"60",
						   33460 => x"00",		-- 0082b4: 0081            
						   33461 => x"81",
						   33462 => x"3C",		-- 0082b6: 3C49             MOV.W   @R9+,R12
						   33463 => x"69",
						   33464 => x"7F",		-- 0082b8: 7F4C             MOV.B   @R12+,R15
						   33465 => x"6C",
						   33466 => x"0F",		-- 0082ba: 0F5F             RLA.W   R15
						   33467 => x"7F",
						   33468 => x"1F",		-- 0082bc: 1F4F             MOV.W   0x80fc(R15),R15
						   33469 => x"6F",
						   33470 => x"FC",		-- 0082be: FC80            
						   33471 => x"80",
						   33472 => x"3D",		-- 0082c0: 3D49             MOV.W   @R9+,R13
						   33473 => x"69",
						   33474 => x"8F",		-- 0082c2: 8F12             CALL    R15
						   33475 => x"32",
						   33476 => x"1A",		-- 0082c4: 1A83             DEC.W   R10
						   33477 => x"A3",
						   33478 => x"F7",		-- 0082c6: F723             JNE     ($C$L21)
						   33479 => x"43",
						   33480 => x"B0",		-- 0082c8: B012             CALL    #_system_post_cinit
						   33481 => x"32",
						   33482 => x"68",		-- 0082ca: 6883            
						   33483 => x"83",
						   33484 => x"30",		-- 0082cc: 3040             BR      #__mspabi_func_epilog_2
						   33485 => x"60",
						   33486 => x"58",		-- 0082ce: 5883            
						   33487 => x"83",
						   -- Begin: __mspabi_slli
						   33488 => x"3D",		-- 0082d0: 3DF0             AND.W   #0x000f,R13
						   33489 => x"10",
						   33490 => x"0F",		-- 0082d2: 0F00            
						   33491 => x"00",
						   33492 => x"3D",		-- 0082d4: 3DE0             XOR.W   #0x000f,R13
						   33493 => x"00",
						   33494 => x"0F",		-- 0082d6: 0F00            
						   33495 => x"00",
						   33496 => x"0D",		-- 0082d8: 0D5D             RLA.W   R13
						   33497 => x"7D",
						   33498 => x"00",		-- 0082da: 005D             ADD.W   R13,PC
						   33499 => x"7D",
						   -- Begin: __mspabi_slli_15
						   33500 => x"0C",		-- 0082dc: 0C5C             RLA.W   R12
						   33501 => x"7C",
						   -- Begin: __mspabi_slli_14
						   33502 => x"0C",		-- 0082de: 0C5C             RLA.W   R12
						   33503 => x"7C",
						   -- Begin: __mspabi_slli_13
						   33504 => x"0C",		-- 0082e0: 0C5C             RLA.W   R12
						   33505 => x"7C",
						   -- Begin: __mspabi_slli_12
						   33506 => x"0C",		-- 0082e2: 0C5C             RLA.W   R12
						   33507 => x"7C",
						   -- Begin: __mspabi_slli_11
						   33508 => x"0C",		-- 0082e4: 0C5C             RLA.W   R12
						   33509 => x"7C",
						   -- Begin: __mspabi_slli_10
						   33510 => x"0C",		-- 0082e6: 0C5C             RLA.W   R12
						   33511 => x"7C",
						   -- Begin: __mspabi_slli_9
						   33512 => x"0C",		-- 0082e8: 0C5C             RLA.W   R12
						   33513 => x"7C",
						   -- Begin: __mspabi_slli_8
						   33514 => x"0C",		-- 0082ea: 0C5C             RLA.W   R12
						   33515 => x"7C",
						   -- Begin: __mspabi_slli_7
						   33516 => x"0C",		-- 0082ec: 0C5C             RLA.W   R12
						   33517 => x"7C",
						   -- Begin: __mspabi_slli_6
						   33518 => x"0C",		-- 0082ee: 0C5C             RLA.W   R12
						   33519 => x"7C",
						   -- Begin: __mspabi_slli_5
						   33520 => x"0C",		-- 0082f0: 0C5C             RLA.W   R12
						   33521 => x"7C",
						   -- Begin: __mspabi_slli_4
						   33522 => x"0C",		-- 0082f2: 0C5C             RLA.W   R12
						   33523 => x"7C",
						   -- Begin: __mspabi_slli_3
						   33524 => x"0C",		-- 0082f4: 0C5C             RLA.W   R12
						   33525 => x"7C",
						   -- Begin: __mspabi_slli_2
						   33526 => x"0C",		-- 0082f6: 0C5C             RLA.W   R12
						   33527 => x"7C",
						   -- Begin: __mspabi_slli_1
						   33528 => x"0C",		-- 0082f8: 0C5C             RLA.W   R12
						   33529 => x"7C",
						   33530 => x"30",		-- 0082fa: 3041             RET     
						   33531 => x"61",
						   -- Begin: _c_int00_noargs
						   33532 => x"31",		-- 0082fc: 3140             MOV.W   #0x3000,SP
						   33533 => x"60",
						   33534 => x"00",		-- 0082fe: 0030            
						   33535 => x"30",
						   33536 => x"B0",		-- 008300: B012             CALL    #_system_pre_init
						   33537 => x"32",
						   33538 => x"64",		-- 008302: 6483            
						   33539 => x"83",
						   33540 => x"0C",		-- 008304: 0C93             TST.W   R12
						   33541 => x"B3",
						   33542 => x"02",		-- 008306: 0224             JEQ     ($C$L2)
						   33543 => x"44",
						   33544 => x"B0",		-- 008308: B012             CALL    #__TI_auto_init_nobinit_nopinit
						   33545 => x"32",
						   33546 => x"8E",		-- 00830a: 8E82            
						   33547 => x"82",
						   33548 => x"0C",		-- 00830c: 0C43             CLR.W   R12
						   33549 => x"63",
						   33550 => x"B0",		-- 00830e: B012             CALL    #main
						   33551 => x"32",
						   33552 => x"04",		-- 008310: 0481            
						   33553 => x"81",
						   33554 => x"1C",		-- 008312: 1C43             MOV.W   #1,R12
						   33555 => x"63",
						   33556 => x"B0",		-- 008314: B012             CALL    #abort
						   33557 => x"32",
						   33558 => x"5E",		-- 008316: 5E83            
						   33559 => x"83",
						   -- Begin: Timer_ISR
						   33560 => x"92",		-- 008318: 9252             ADD.W   &frequency,&TB0CCR0_L
						   33561 => x"72",
						   33562 => x"00",		-- 00831a: 0021            
						   33563 => x"21",
						   33564 => x"92",		-- 00831c: 9203            
						   33565 => x"03",
						   33566 => x"F2",		-- 00831e: F2E0             XOR.B   #0x0010,&P2OUT
						   33567 => x"00",
						   33568 => x"10",		-- 008320: 1000            
						   33569 => x"00",
						   33570 => x"03",		-- 008322: 0302            
						   33571 => x"02",
						   33572 => x"92",		-- 008324: 92C3             BIC.W   #1,&TB0CCTL0_L
						   33573 => x"E3",
						   33574 => x"82",		-- 008326: 8203            
						   33575 => x"03",
						   33576 => x"00",		-- 008328: 0013             RETI    
						   33577 => x"33",
						   -- Begin: __TI_decompress_none
						   33578 => x"0F",		-- 00832a: 0F4C             MOV.W   R12,R15
						   33579 => x"6C",
						   33580 => x"0C",		-- 00832c: 0C4D             MOV.W   R13,R12
						   33581 => x"6D",
						   33582 => x"3D",		-- 00832e: 3D40             MOV.W   #0x0003,R13
						   33583 => x"60",
						   33584 => x"03",		-- 008330: 0300            
						   33585 => x"00",
						   33586 => x"0D",		-- 008332: 0D5F             ADD.W   R15,R13
						   33587 => x"7F",
						   33588 => x"1E",		-- 008334: 1E4F             MOV.W   0x0001(R15),R14
						   33589 => x"6F",
						   33590 => x"01",		-- 008336: 0100            
						   33591 => x"00",
						   33592 => x"30",		-- 008338: 3040             BR      #memcpy
						   33593 => x"60",
						   33594 => x"3C",		-- 00833a: 3C83            
						   33595 => x"83",
						   -- Begin: memcpy
						   33596 => x"0E",		-- 00833c: 0E93             TST.W   R14
						   33597 => x"B3",
						   33598 => x"06",		-- 00833e: 0624             JEQ     ($C$L2)
						   33599 => x"44",
						   33600 => x"0F",		-- 008340: 0F4C             MOV.W   R12,R15
						   33601 => x"6C",
						   33602 => x"1F",		-- 008342: 1F53             INC.W   R15
						   33603 => x"73",
						   33604 => x"FF",		-- 008344: FF4D             MOV.B   @R13+,0xffff(R15)
						   33605 => x"6D",
						   33606 => x"FF",		-- 008346: FFFF            
						   33607 => x"FF",
						   33608 => x"1E",		-- 008348: 1E83             DEC.W   R14
						   33609 => x"A3",
						   33610 => x"FB",		-- 00834a: FB23             JNE     ($C$L1)
						   33611 => x"43",
						   33612 => x"30",		-- 00834c: 3041             RET     
						   33613 => x"61",
						   -- Begin: __mspabi_func_epilog_7
						   -- Begin: __mspabi_func_epilog
						   33614 => x"34",		-- 00834e: 3441             POP.W   R4
						   33615 => x"61",
						   -- Begin: __mspabi_func_epilog_6
						   33616 => x"35",		-- 008350: 3541             POP.W   R5
						   33617 => x"61",
						   -- Begin: __mspabi_func_epilog_5
						   33618 => x"36",		-- 008352: 3641             POP.W   R6
						   33619 => x"61",
						   -- Begin: __mspabi_func_epilog_4
						   33620 => x"37",		-- 008354: 3741             POP.W   R7
						   33621 => x"61",
						   -- Begin: __mspabi_func_epilog_3
						   33622 => x"38",		-- 008356: 3841             POP.W   R8
						   33623 => x"61",
						   -- Begin: __mspabi_func_epilog_2
						   33624 => x"39",		-- 008358: 3941             POP.W   R9
						   33625 => x"61",
						   -- Begin: __mspabi_func_epilog_1
						   33626 => x"3A",		-- 00835a: 3A41             POP.W   R10
						   33627 => x"61",
						   33628 => x"30",		-- 00835c: 3041             RET     
						   33629 => x"61",
						   -- Begin: abort
						   33630 => x"03",		-- 00835e: 0343             NOP     
						   33631 => x"63",
						   33632 => x"FF",		-- 008360: FF3F             JMP     ($C$L1)
						   33633 => x"5F",
						   33634 => x"03",		-- 008362: 0343             NOP     
						   33635 => x"63",
						   -- Begin: _system_pre_init
						   33636 => x"1C",		-- 008364: 1C43             MOV.W   #1,R12
						   33637 => x"63",
						   33638 => x"30",		-- 008366: 3041             RET     
						   33639 => x"61",
						   -- Begin: _system_post_cinit
						   33640 => x"30",		-- 008368: 3041             RET     
						   33641 => x"61",
						   -- ISR Trap
						   33642 => x"32",		-- 00836a: 32D0             BIS.W   #0x0010,SR
						   33643 => x"F0",
						   33644 => x"10",		-- 00836c: 1000            
						   33645 => x"00",
						   33646 => x"FD",		-- 00836e: FD3F             JMP     (__TI_ISR_TRAP)
						   33647 => x"5F",
						   33648 => x"03",		-- 008370: 0343             NOP     
						   33649 => x"63",
						   -- IRQ Vectors (Interrupt Vectors)
						   65486 => x"6a",		-- 00ffce:836a PORT4 __TI_int22 int22
						   65487 => x"83",
						   65488 => x"6a",		-- 00ffd0:836a PORT3 __TI_int23 int23
						   65489 => x"83",
						   65490 => x"6a",		-- 00ffd2:836a PORT2 __TI_int24 int24
						   65491 => x"83",
						   65492 => x"6a",		-- 00ffd4:836a PORT1 __TI_int25 int25
						   65493 => x"83",
						   65494 => x"6a",		-- 00ffd6:836a SAC1_SAC3 __TI_int26 int26
						   65495 => x"83",
						   65496 => x"6a",		-- 00ffd8:836a SAC0_SAC2 __TI_int27 int27
						   65497 => x"83",
						   65498 => x"6a",		-- 00ffda:836a ECOMP0_ECOMP1 __TI_int28 int28
						   65499 => x"83",
						   65500 => x"6a",		-- 00ffdc:836a ADC __TI_int29 int29
						   65501 => x"83",
						   65502 => x"6a",		-- 00ffde:836a EUSCI_B1 __TI_int30 int30
						   65503 => x"83",
						   65504 => x"6a",		-- 00ffe0:836a EUSCI_B0 __TI_int31 int31
						   65505 => x"83",
						   65506 => x"6a",		-- 00ffe2:836a EUSCI_A1 __TI_int32 int32
						   65507 => x"83",
						   65508 => x"6a",		-- 00ffe4:836a EUSCI_A0 __TI_int33 int33
						   65509 => x"83",
						   65510 => x"6a",		-- 00ffe6:836a WDT __TI_int34 int34
						   65511 => x"83",
						   65512 => x"6a",		-- 00ffe8:836a RTC __TI_int35 int35
						   65513 => x"83",
						   65514 => x"6a",		-- 00ffea:836a TIMER3_B1 __TI_int36 int36
						   65515 => x"83",
						   65516 => x"6a",		-- 00ffec:836a TIMER3_B0 __TI_int37 int37
						   65517 => x"83",
						   65518 => x"6a",		-- 00ffee:836a TIMER2_B1 __TI_int38 int38
						   65519 => x"83",
						   65520 => x"6a",		-- 00fff0:836a TIMER2_B0 __TI_int39 int39
						   65521 => x"83",
						   65522 => x"6a",		-- 00fff2:836a TIMER1_B1 __TI_int40 int40
						   65523 => x"83",
						   65524 => x"6a",		-- 00fff4:836a TIMER1_B0 __TI_int41 int41
						   65525 => x"83",
						   65526 => x"6a",		-- 00fff6:836a TIMER0_B1 __TI_int42 int42
						   65527 => x"83",
						   65528 => x"18",		-- 00fff8:8318 TIMER0_B0 __TI_int43 int43
						   65529 => x"83",
						   65530 => x"6a",		-- 00fffa:836a UNMI __TI_int44 int44
						   65531 => x"83",
						   65532 => x"6a",		-- 00fffc:836a SYSNMI __TI_int45 int45
						   65533 => x"83",
						   65534 => x"fc",		-- 00fffe:82fc .reset _reset_vector reset
						   65535 => x"82",
						   others => x"00");

    signal EN : std_logic;
    
    begin
    -- Note 1:  The bus system uses a 16-bit Address (MAB)
    --          This address size can access locations from x0000 to xFFFF
    --          But our array is only defined from x8000 to xFFFF and
    --          if we try to access it with any other address, it will crash.
    --          So the first thing we need to do is create a local enable that
    --          will only assert when MAB is within x8000 to xFFFF.

     LOCAL_EN : process (MAB) 
     begin
         if ( (to_integer(unsigned(MAB)) >= 32768) and (to_integer(unsigned(MAB)) <= 65535)) then
           EN <= '1';
         else 
           EN <= '0';
         end if;
     end process;

    
    -- Note 2:  The bus system uses a 16-bit Address (MAB)
    --          The MDB_out is also provided as a 16-bit word
    --          However, the memory array is actually built as 8-bit bytes.
    --          So for a given 16-bit MAB, we give MDB_out = HB : LB
    --                                                 or  = ROM(MAB);1) : ROM(MAB)

    MEMORY_ROM : process (clk) 
    begin
        if (rising_edge(clk)) then
            if (EN='1' and write='0') then
                if(Byte = '0') then                      
                    MDB_in <= ROM(to_integer(unsigned(MAB)) + 1 ) & ROM(to_integer(unsigned(MAB)));
                else
                    MDB_in <= x"00" & ROM(to_integer(unsigned(MAB)));
                end if;
            end if;
        end if;
    end process;


end architecture;