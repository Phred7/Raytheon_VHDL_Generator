library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;


entity highroller_memory is
    port ( clk	: in	std_logic;
         MAB		: in	std_logic_vector(15 downto 0);
         MDB_in  	: out	std_logic_vector(15 downto 0);
         MDB_out  	: in	std_logic_vector(15 downto 0);
         write	    : in	std_logic;
         Byte       : in    std_logic);
end entity;

architecture highroller_memory_arch of highroller_memory is

type rom_type is array (32768 to 65535) of std_logic_vector(7 downto 0);  -- this is MAB: x8000 to xFFFF
    
constant ROM : rom_type :=(						   33792 => x"02",
						   33793 => x"00",
						   33794 => x"fe",
						   33795 => x"00",
						   33806 => x"12",
						   33807 => x"00",
						   33808 => x"01",
						   33809 => x"00",
						   33818 => x"22",
						   33819 => x"00",
						   33820 => x"02",
						   33821 => x"00",
						   33830 => x"24",
						   33831 => x"00",
						   33926 => x"02",
						   33927 => x"00",
						   33928 => x"4e",
						   33929 => x"d6",
						   33930 => x"aa",
						   33931 => x"da",
						   33932 => x"78",
						   33933 => x"d7",
						   33934 => x"b4",
						   33935 => x"d6",
						   33936 => x"ac",
						   33937 => x"d1",
						   33938 => x"b8",
						   33939 => x"db",
						   33940 => x"7c",
						   33941 => x"d5",
						   33994 => x"78",
						   33995 => x"20",
						   33998 => x"78",
						   33999 => x"20",
						   34000 => x"01",
						   34001 => x"00",
						   34002 => x"78",
						   34003 => x"20",
						   34004 => x"02",
						   34005 => x"00",
						   34038 => x"dc",
						   34039 => x"e1",
						   34040 => x"dc",
						   34041 => x"e1",
						   34042 => x"03",
						   34043 => x"00",
						   34046 => x"01",
						   34047 => x"00",
						   34050 => x"c4",
						   34051 => x"e0",
						   34052 => x"b8",
						   34053 => x"d2",
						   34054 => x"3a",
						   34055 => x"e1",
						   34058 => x"aa",
						   34059 => x"00",
						   34060 => x"00",
						   34061 => x"84",
						   34062 => x"00",
						   34063 => x"20",
						   34064 => x"08",
						   34065 => x"85",
						   34066 => x"fe",
						   34067 => x"20",
						   -- Begin: program memory TEXT Section
						   56500 => x"31",		-- 00dcb4: 3182             SUB.W   #8,SP
						   56501 => x"A2",
						   56502 => x"B2",		-- 00dcb6: B240             MOV.W   #0x5a80,&WDTCTL_L
						   56503 => x"60",
						   56504 => x"80",		-- 00dcb8: 805A            
						   56505 => x"5A",
						   56506 => x"CC",		-- 00dcba: CC01            
						   56507 => x"01",
						   56508 => x"81",		-- 00dcbc: 8143             CLR.W   0x0004(SP)
						   56509 => x"63",
						   56510 => x"04",		-- 00dcbe: 0400            
						   56511 => x"00",
						   56512 => x"1C",		-- 00dcc0: 1C41             MOV.W   0x0002(SP),R12
						   56513 => x"61",
						   56514 => x"02",		-- 00dcc2: 0200            
						   56515 => x"00",
						   56516 => x"B0",		-- 00dcc4: B012             CALL    #buff_value
						   56517 => x"32",
						   56518 => x"28",		-- 00dcc6: 28E1            
						   56519 => x"E1",
						   56520 => x"1C",		-- 00dcc8: 1C41             MOV.W   0x0006(SP),R12
						   56521 => x"61",
						   56522 => x"06",		-- 00dcca: 0600            
						   56523 => x"00",
						   56524 => x"B0",		-- 00dccc: B012             CALL    #buff_value
						   56525 => x"32",
						   56526 => x"28",		-- 00dcce: 28E1            
						   56527 => x"E1",
						   56528 => x"81",		-- 00dcd0: 8193             TST.W   0x0004(SP)
						   56529 => x"B3",
						   56530 => x"04",		-- 00dcd2: 0400            
						   56531 => x"00",
						   56532 => x"06",		-- 00dcd4: 0620             JNE     ($C$L1)
						   56533 => x"40",
						   56534 => x"B1",		-- 00dcd6: B140             MOV.W   #0x852c,0x0000(SP)
						   56535 => x"60",
						   56536 => x"2C",		-- 00dcd8: 2C85            
						   56537 => x"85",
						   56538 => x"00",		-- 00dcda: 0000            
						   56539 => x"00",
						   56540 => x"B0",		-- 00dcdc: B012             CALL    #printf
						   56541 => x"32",
						   56542 => x"F2",		-- 00dcde: F2DC            
						   56543 => x"DC",
						   56544 => x"05",		-- 00dce0: 053C             JMP     ($C$L2)
						   56545 => x"5C",
						   56546 => x"B1",		-- 00dce2: B140             MOV.W   #0x852c,0x0000(SP)
						   56547 => x"60",
						   56548 => x"2C",		-- 00dce4: 2C85            
						   56549 => x"85",
						   56550 => x"00",		-- 00dce6: 0000            
						   56551 => x"00",
						   56552 => x"B0",		-- 00dce8: B012             CALL    #printf
						   56553 => x"32",
						   56554 => x"F2",		-- 00dcea: F2DC            
						   56555 => x"DC",
						   56556 => x"0C",		-- 00dcec: 0C43             CLR.W   R12
						   56557 => x"63",
						   56558 => x"31",		-- 00dcee: 3152             ADD.W   #8,SP
						   56559 => x"72",
						   56560 => x"30",		-- 00dcf0: 3041             RET     
						   56561 => x"61",
						   -- Begin: printf
						   56562 => x"0A",		-- 00dcf2: 0A12             PUSH    R10
						   56563 => x"32",
						   56564 => x"21",		-- 00dcf4: 2183             DECD.W  SP
						   56565 => x"A3",
						   56566 => x"92",		-- 00dcf6: 9212             CALL    &_lock
						   56567 => x"32",
						   56568 => x"F2",		-- 00dcf8: F220            
						   56569 => x"20",
						   56570 => x"B2",		-- 00dcfa: B293             CMP.W   #-1,&0x200c
						   56571 => x"B3",
						   56572 => x"0C",		-- 00dcfc: 0C20            
						   56573 => x"20",
						   56574 => x"02",		-- 00dcfe: 0220             JNE     ($C$L1)
						   56575 => x"40",
						   56576 => x"3A",		-- 00dd00: 3A43             MOV.W   #-1,R10
						   56577 => x"63",
						   56578 => x"0F",		-- 00dd02: 0F3C             JMP     ($C$L2)
						   56579 => x"5C",
						   56580 => x"B1",		-- 00dd04: B140             MOV.W   #0xe1d4,0x0000(SP)
						   56581 => x"60",
						   56582 => x"D4",		-- 00dd06: D4E1            
						   56583 => x"E1",
						   56584 => x"00",		-- 00dd08: 0000            
						   56585 => x"00",
						   56586 => x"0D",		-- 00dd0a: 0D41             MOV.W   SP,R13
						   56587 => x"61",
						   56588 => x"3D",		-- 00dd0c: 3D52             ADD.W   #8,R13
						   56589 => x"72",
						   56590 => x"3E",		-- 00dd0e: 3E40             MOV.W   #0x200c,R14
						   56591 => x"60",
						   56592 => x"0C",		-- 00dd10: 0C20            
						   56593 => x"20",
						   56594 => x"0C",		-- 00dd12: 0C41             MOV.W   SP,R12
						   56595 => x"61",
						   56596 => x"3C",		-- 00dd14: 3C50             ADD.W   #0x0006,R12
						   56597 => x"70",
						   56598 => x"06",		-- 00dd16: 0600            
						   56599 => x"00",
						   56600 => x"3F",		-- 00dd18: 3F40             MOV.W   #0xe1c8,R15
						   56601 => x"60",
						   56602 => x"C8",		-- 00dd1a: C8E1            
						   56603 => x"E1",
						   56604 => x"B0",		-- 00dd1c: B012             CALL    #__TI_printfi
						   56605 => x"32",
						   56606 => x"24",		-- 00dd1e: 24AC            
						   56607 => x"AC",
						   56608 => x"0A",		-- 00dd20: 0A4C             MOV.W   R12,R10
						   56609 => x"6C",
						   56610 => x"92",		-- 00dd22: 9212             CALL    &_unlock
						   56611 => x"32",
						   56612 => x"F4",		-- 00dd24: F420            
						   56613 => x"20",
						   56614 => x"0C",		-- 00dd26: 0C4A             MOV.W   R10,R12
						   56615 => x"6A",
						   56616 => x"21",		-- 00dd28: 2153             INCD.W  SP
						   56617 => x"73",
						   56618 => x"3A",		-- 00dd2a: 3A41             POP.W   R10
						   56619 => x"61",
						   56620 => x"30",		-- 00dd2c: 3041             RET     
						   56621 => x"61",
						   -- Begin: __TI_cleanup
						   56622 => x"0A",		-- 00dd2e: 0A12             PUSH    R10
						   56623 => x"32",
						   56624 => x"09",		-- 00dd30: 0912             PUSH    R9
						   56625 => x"32",
						   56626 => x"3C",		-- 00dd32: 3C40             MOV.W   #0x2000,R12
						   56627 => x"60",
						   56628 => x"00",		-- 00dd34: 0020            
						   56629 => x"20",
						   56630 => x"B0",		-- 00dd36: B012             CALL    #__TI_closefile
						   56631 => x"32",
						   56632 => x"28",		-- 00dd38: 28D4            
						   56633 => x"D4",
						   56634 => x"A2",		-- 00dd3a: A293             CMP.W   #2,&__TI_ft_end
						   56635 => x"B3",
						   56636 => x"F6",		-- 00dd3c: F620            
						   56637 => x"20",
						   56638 => x"0F",		-- 00dd3e: 0F38             JL      ($C$L37)
						   56639 => x"58",
						   56640 => x"3A",		-- 00dd40: 3A40             MOV.W   #0x200c,R10
						   56641 => x"60",
						   56642 => x"0C",		-- 00dd42: 0C20            
						   56643 => x"20",
						   56644 => x"19",		-- 00dd44: 1943             MOV.W   #1,R9
						   56645 => x"63",
						   56646 => x"8A",		-- 00dd46: 8A93             TST.W   0x0000(R10)
						   56647 => x"B3",
						   56648 => x"00",		-- 00dd48: 0000            
						   56649 => x"00",
						   56650 => x"03",		-- 00dd4a: 0338             JL      ($C$L36)
						   56651 => x"58",
						   56652 => x"0C",		-- 00dd4c: 0C4A             MOV.W   R10,R12
						   56653 => x"6A",
						   56654 => x"B0",		-- 00dd4e: B012             CALL    #__TI_closefile
						   56655 => x"32",
						   56656 => x"28",		-- 00dd50: 28D4            
						   56657 => x"D4",
						   56658 => x"3A",		-- 00dd52: 3A50             ADD.W   #0x000c,R10
						   56659 => x"70",
						   56660 => x"0C",		-- 00dd54: 0C00            
						   56661 => x"00",
						   56662 => x"19",		-- 00dd56: 1953             INC.W   R9
						   56663 => x"73",
						   56664 => x"19",		-- 00dd58: 1992             CMP.W   &__TI_ft_end,R9
						   56665 => x"B2",
						   56666 => x"F6",		-- 00dd5a: F620            
						   56667 => x"20",
						   56668 => x"F4",		-- 00dd5c: F43B             JL      ($C$L35)
						   56669 => x"5B",
						   56670 => x"30",		-- 00dd5e: 3040             BR      #__mspabi_func_epilog_2
						   56671 => x"60",
						   56672 => x"7A",		-- 00dd60: 7AE1            
						   56673 => x"E1",
						   -- Begin: finddevice
						   56674 => x"0A",		-- 00dd62: 0A12             PUSH    R10
						   56675 => x"32",
						   56676 => x"09",		-- 00dd64: 0912             PUSH    R9
						   56677 => x"32",
						   56678 => x"08",		-- 00dd66: 0812             PUSH    R8
						   56679 => x"32",
						   56680 => x"08",		-- 00dd68: 084C             MOV.W   R12,R8
						   56681 => x"6C",
						   56682 => x"C8",		-- 00dd6a: C893             TST.B   0x0000(R8)
						   56683 => x"B3",
						   56684 => x"00",		-- 00dd6c: 0000            
						   56685 => x"00",
						   56686 => x"10",		-- 00dd6e: 1024             JEQ     ($C$L3)
						   56687 => x"44",
						   56688 => x"3A",		-- 00dd70: 3A40             MOV.W   #0x2092,R10
						   56689 => x"60",
						   56690 => x"92",		-- 00dd72: 9220            
						   56691 => x"20",
						   56692 => x"29",		-- 00dd74: 2943             MOV.W   #2,R9
						   56693 => x"63",
						   56694 => x"0C",		-- 00dd76: 0C4A             MOV.W   R10,R12
						   56695 => x"6A",
						   56696 => x"0D",		-- 00dd78: 0D48             MOV.W   R8,R13
						   56697 => x"68",
						   56698 => x"B0",		-- 00dd7a: B012             CALL    #strcmp
						   56699 => x"32",
						   56700 => x"96",		-- 00dd7c: 96E0            
						   56701 => x"E0",
						   56702 => x"0C",		-- 00dd7e: 0C93             TST.W   R12
						   56703 => x"B3",
						   56704 => x"03",		-- 00dd80: 0320             JNE     ($C$L2)
						   56705 => x"40",
						   56706 => x"0C",		-- 00dd82: 0C4A             MOV.W   R10,R12
						   56707 => x"6A",
						   56708 => x"30",		-- 00dd84: 3040             BR      #__mspabi_func_epilog_3
						   56709 => x"60",
						   56710 => x"78",		-- 00dd86: 78E1            
						   56711 => x"E1",
						   56712 => x"3A",		-- 00dd88: 3A50             ADD.W   #0x001a,R10
						   56713 => x"70",
						   56714 => x"1A",		-- 00dd8a: 1A00            
						   56715 => x"00",
						   56716 => x"19",		-- 00dd8c: 1983             DEC.W   R9
						   56717 => x"A3",
						   56718 => x"F3",		-- 00dd8e: F323             JNE     ($C$L1)
						   56719 => x"43",
						   56720 => x"0C",		-- 00dd90: 0C43             CLR.W   R12
						   56721 => x"63",
						   56722 => x"30",		-- 00dd92: 3040             BR      #__mspabi_func_epilog_3
						   56723 => x"60",
						   56724 => x"78",		-- 00dd94: 78E1            
						   56725 => x"E1",
						   -- Begin: __TI_writemsg
						   56726 => x"82",		-- 00dd96: 824F             MOV.W   R15,&_CIOBUF_
						   56727 => x"6F",
						   56728 => x"00",		-- 00dd98: 0080            
						   56729 => x"80",
						   56730 => x"C2",		-- 00dd9a: C24C             MOV.B   R12,&0x8002
						   56731 => x"6C",
						   56732 => x"02",		-- 00dd9c: 0280            
						   56733 => x"80",
						   56734 => x"3C",		-- 00dd9e: 3C40             MOV.W   #0x8003,R12
						   56735 => x"60",
						   56736 => x"03",		-- 00dda0: 0380            
						   56737 => x"80",
						   56738 => x"3B",		-- 00dda2: 3B42             MOV.W   #8,R11
						   56739 => x"62",
						   56740 => x"1C",		-- 00dda4: 1C53             INC.W   R12
						   56741 => x"73",
						   56742 => x"FC",		-- 00dda6: FC4D             MOV.B   @R13+,0xffff(R12)
						   56743 => x"6D",
						   56744 => x"FF",		-- 00dda8: FFFF            
						   56745 => x"FF",
						   56746 => x"1B",		-- 00ddaa: 1B83             DEC.W   R11
						   56747 => x"A3",
						   56748 => x"FB",		-- 00ddac: FB23             JNE     ($C$L1)
						   56749 => x"43",
						   56750 => x"0F",		-- 00ddae: 0F93             TST.W   R15
						   56751 => x"B3",
						   56752 => x"07",		-- 00ddb0: 0724             JEQ     (C$$IO$$)
						   56753 => x"44",
						   56754 => x"3D",		-- 00ddb2: 3D40             MOV.W   #0x800b,R13
						   56755 => x"60",
						   56756 => x"0B",		-- 00ddb4: 0B80            
						   56757 => x"80",
						   56758 => x"1D",		-- 00ddb6: 1D53             INC.W   R13
						   56759 => x"73",
						   56760 => x"FD",		-- 00ddb8: FD4E             MOV.B   @R14+,0xffff(R13)
						   56761 => x"6E",
						   56762 => x"FF",		-- 00ddba: FFFF            
						   56763 => x"FF",
						   56764 => x"1F",		-- 00ddbc: 1F83             DEC.W   R15
						   56765 => x"A3",
						   56766 => x"FB",		-- 00ddbe: FB23             JNE     ($C$L2)
						   56767 => x"43",
						   56768 => x"03",		-- 00ddc0: 0343             NOP     
						   56769 => x"63",
						   56770 => x"30",		-- 00ddc2: 3041             RET     
						   56771 => x"61",
						   -- Begin: __mspabi_subd
						   56772 => x"31",		-- 00ddc4: 3182             SUB.W   #8,SP
						   56773 => x"A2",
						   56774 => x"81",		-- 00ddc6: 814C             MOV.W   R12,0x0000(SP)
						   56775 => x"6C",
						   56776 => x"00",		-- 00ddc8: 0000            
						   56777 => x"00",
						   56778 => x"81",		-- 00ddca: 814D             MOV.W   R13,0x0002(SP)
						   56779 => x"6D",
						   56780 => x"02",		-- 00ddcc: 0200            
						   56781 => x"00",
						   56782 => x"81",		-- 00ddce: 814E             MOV.W   R14,0x0004(SP)
						   56783 => x"6E",
						   56784 => x"04",		-- 00ddd0: 0400            
						   56785 => x"00",
						   56786 => x"81",		-- 00ddd2: 814F             MOV.W   R15,0x0006(SP)
						   56787 => x"6F",
						   56788 => x"06",		-- 00ddd4: 0600            
						   56789 => x"00",
						   56790 => x"F1",		-- 00ddd6: F1E0             XOR.B   #0x0080,0x0007(SP)
						   56791 => x"00",
						   56792 => x"80",		-- 00ddd8: 8000            
						   56793 => x"00",
						   56794 => x"07",		-- 00ddda: 0700            
						   56795 => x"00",
						   56796 => x"2C",		-- 00dddc: 2C41             MOV.W   @SP,R12
						   56797 => x"61",
						   56798 => x"1D",		-- 00ddde: 1D41             MOV.W   0x0002(SP),R13
						   56799 => x"61",
						   56800 => x"02",		-- 00dde0: 0200            
						   56801 => x"00",
						   56802 => x"1E",		-- 00dde2: 1E41             MOV.W   0x0004(SP),R14
						   56803 => x"61",
						   56804 => x"04",		-- 00dde4: 0400            
						   56805 => x"00",
						   56806 => x"1F",		-- 00dde6: 1F41             MOV.W   0x0006(SP),R15
						   56807 => x"61",
						   56808 => x"06",		-- 00dde8: 0600            
						   56809 => x"00",
						   56810 => x"B0",		-- 00ddea: B012             CALL    #__mspabi_addd
						   56811 => x"32",
						   56812 => x"56",		-- 00ddec: 569A            
						   56813 => x"9A",
						   56814 => x"31",		-- 00ddee: 3152             ADD.W   #8,SP
						   56815 => x"72",
						   56816 => x"30",		-- 00ddf0: 3041             RET     
						   56817 => x"61",
						   -- Begin: copysignl
						   -- Begin: copysign
						   56818 => x"0A",		-- 00ddf2: 0A12             PUSH    R10
						   56819 => x"32",
						   56820 => x"1A",		-- 00ddf4: 1A41             MOV.W   0x0008(SP),R10
						   56821 => x"61",
						   56822 => x"08",		-- 00ddf6: 0800            
						   56823 => x"00",
						   56824 => x"1B",		-- 00ddf8: 1B41             MOV.W   0x000a(SP),R11
						   56825 => x"61",
						   56826 => x"0A",		-- 00ddfa: 0A00            
						   56827 => x"00",
						   56828 => x"0A",		-- 00ddfc: 0AF3             AND.W   #0,R10
						   56829 => x"13",
						   56830 => x"3B",		-- 00ddfe: 3BF0             AND.W   #0x8000,R11
						   56831 => x"10",
						   56832 => x"00",		-- 00de00: 0080            
						   56833 => x"80",
						   56834 => x"3E",		-- 00de02: 3EF3             AND.W   #-1,R14
						   56835 => x"13",
						   56836 => x"3F",		-- 00de04: 3FF0             AND.W   #0x7fff,R15
						   56837 => x"10",
						   56838 => x"FF",		-- 00de06: FF7F            
						   56839 => x"7F",
						   56840 => x"0E",		-- 00de08: 0EDA             BIS.W   R10,R14
						   56841 => x"FA",
						   56842 => x"0F",		-- 00de0a: 0FDB             BIS.W   R11,R15
						   56843 => x"FB",
						   56844 => x"0B",		-- 00de0c: 0B43             CLR.W   R11
						   56845 => x"63",
						   56846 => x"0B",		-- 00de0e: 0BDD             BIS.W   R13,R11
						   56847 => x"FD",
						   56848 => x"0D",		-- 00de10: 0D43             CLR.W   R13
						   56849 => x"63",
						   56850 => x"0D",		-- 00de12: 0DDC             BIS.W   R12,R13
						   56851 => x"FC",
						   56852 => x"0E",		-- 00de14: 0ED3             BIS.W   #0,R14
						   56853 => x"F3",
						   56854 => x"0F",		-- 00de16: 0FD3             BIS.W   #0,R15
						   56855 => x"F3",
						   56856 => x"0C",		-- 00de18: 0C4D             MOV.W   R13,R12
						   56857 => x"6D",
						   56858 => x"0D",		-- 00de1a: 0D4B             MOV.W   R11,R13
						   56859 => x"6B",
						   56860 => x"3A",		-- 00de1c: 3A41             POP.W   R10
						   56861 => x"61",
						   56862 => x"30",		-- 00de1e: 3041             RET     
						   56863 => x"61",
						   -- Begin: __TI_readmsg
						   56864 => x"1F",		-- 00de20: 1F42             MOV.W   &_CIOBUF_,R15
						   56865 => x"62",
						   56866 => x"00",		-- 00de22: 0080            
						   56867 => x"80",
						   56868 => x"3B",		-- 00de24: 3B40             MOV.W   #0x8002,R11
						   56869 => x"60",
						   56870 => x"02",		-- 00de26: 0280            
						   56871 => x"80",
						   56872 => x"3E",		-- 00de28: 3E42             MOV.W   #8,R14
						   56873 => x"62",
						   56874 => x"1C",		-- 00de2a: 1C53             INC.W   R12
						   56875 => x"73",
						   56876 => x"FC",		-- 00de2c: FC4B             MOV.B   @R11+,0xffff(R12)
						   56877 => x"6B",
						   56878 => x"FF",		-- 00de2e: FFFF            
						   56879 => x"FF",
						   56880 => x"1E",		-- 00de30: 1E83             DEC.W   R14
						   56881 => x"A3",
						   56882 => x"FB",		-- 00de32: FB23             JNE     ($C$L4)
						   56883 => x"43",
						   56884 => x"0D",		-- 00de34: 0D93             TST.W   R13
						   56885 => x"B3",
						   56886 => x"09",		-- 00de36: 0924             JEQ     ($C$L6)
						   56887 => x"44",
						   56888 => x"0F",		-- 00de38: 0F93             TST.W   R15
						   56889 => x"B3",
						   56890 => x"07",		-- 00de3a: 0724             JEQ     ($C$L6)
						   56891 => x"44",
						   56892 => x"3E",		-- 00de3c: 3E40             MOV.W   #0x800a,R14
						   56893 => x"60",
						   56894 => x"0A",		-- 00de3e: 0A80            
						   56895 => x"80",
						   56896 => x"1D",		-- 00de40: 1D53             INC.W   R13
						   56897 => x"73",
						   56898 => x"FD",		-- 00de42: FD4E             MOV.B   @R14+,0xffff(R13)
						   56899 => x"6E",
						   56900 => x"FF",		-- 00de44: FFFF            
						   56901 => x"FF",
						   56902 => x"1F",		-- 00de46: 1F83             DEC.W   R15
						   56903 => x"A3",
						   56904 => x"FB",		-- 00de48: FB23             JNE     ($C$L5)
						   56905 => x"43",
						   56906 => x"30",		-- 00de4a: 3041             RET     
						   56907 => x"61",
						   -- Begin: __mspabi_srai
						   56908 => x"3D",		-- 00de4c: 3DF0             AND.W   #0x000f,R13
						   56909 => x"10",
						   56910 => x"0F",		-- 00de4e: 0F00            
						   56911 => x"00",
						   56912 => x"3D",		-- 00de50: 3DE0             XOR.W   #0x000f,R13
						   56913 => x"00",
						   56914 => x"0F",		-- 00de52: 0F00            
						   56915 => x"00",
						   56916 => x"0D",		-- 00de54: 0D5D             RLA.W   R13
						   56917 => x"7D",
						   56918 => x"00",		-- 00de56: 005D             ADD.W   R13,PC
						   56919 => x"7D",
						   -- Begin: __mspabi_srai_15
						   56920 => x"0C",		-- 00de58: 0C11             RRA     R12
						   56921 => x"31",
						   -- Begin: __mspabi_srai_14
						   56922 => x"0C",		-- 00de5a: 0C11             RRA     R12
						   56923 => x"31",
						   -- Begin: __mspabi_srai_13
						   56924 => x"0C",		-- 00de5c: 0C11             RRA     R12
						   56925 => x"31",
						   -- Begin: __mspabi_srai_12
						   56926 => x"0C",		-- 00de5e: 0C11             RRA     R12
						   56927 => x"31",
						   -- Begin: __mspabi_srai_11
						   56928 => x"0C",		-- 00de60: 0C11             RRA     R12
						   56929 => x"31",
						   -- Begin: __mspabi_srai_10
						   56930 => x"0C",		-- 00de62: 0C11             RRA     R12
						   56931 => x"31",
						   -- Begin: __mspabi_srai_9
						   56932 => x"0C",		-- 00de64: 0C11             RRA     R12
						   56933 => x"31",
						   -- Begin: __mspabi_srai_8
						   56934 => x"0C",		-- 00de66: 0C11             RRA     R12
						   56935 => x"31",
						   -- Begin: __mspabi_srai_7
						   56936 => x"0C",		-- 00de68: 0C11             RRA     R12
						   56937 => x"31",
						   -- Begin: __mspabi_srai_6
						   56938 => x"0C",		-- 00de6a: 0C11             RRA     R12
						   56939 => x"31",
						   -- Begin: __mspabi_srai_5
						   56940 => x"0C",		-- 00de6c: 0C11             RRA     R12
						   56941 => x"31",
						   -- Begin: __mspabi_srai_4
						   56942 => x"0C",		-- 00de6e: 0C11             RRA     R12
						   56943 => x"31",
						   -- Begin: __mspabi_srai_3
						   56944 => x"0C",		-- 00de70: 0C11             RRA     R12
						   56945 => x"31",
						   -- Begin: __mspabi_srai_2
						   56946 => x"0C",		-- 00de72: 0C11             RRA     R12
						   56947 => x"31",
						   -- Begin: __mspabi_srai_1
						   56948 => x"0C",		-- 00de74: 0C11             RRA     R12
						   56949 => x"31",
						   56950 => x"30",		-- 00de76: 3041             RET     
						   56951 => x"61",
						   -- Begin: __mspabi_slli
						   56952 => x"3D",		-- 00de78: 3DF0             AND.W   #0x000f,R13
						   56953 => x"10",
						   56954 => x"0F",		-- 00de7a: 0F00            
						   56955 => x"00",
						   56956 => x"3D",		-- 00de7c: 3DE0             XOR.W   #0x000f,R13
						   56957 => x"00",
						   56958 => x"0F",		-- 00de7e: 0F00            
						   56959 => x"00",
						   56960 => x"0D",		-- 00de80: 0D5D             RLA.W   R13
						   56961 => x"7D",
						   56962 => x"00",		-- 00de82: 005D             ADD.W   R13,PC
						   56963 => x"7D",
						   -- Begin: __mspabi_slli_15
						   56964 => x"0C",		-- 00de84: 0C5C             RLA.W   R12
						   56965 => x"7C",
						   -- Begin: __mspabi_slli_14
						   56966 => x"0C",		-- 00de86: 0C5C             RLA.W   R12
						   56967 => x"7C",
						   -- Begin: __mspabi_slli_13
						   56968 => x"0C",		-- 00de88: 0C5C             RLA.W   R12
						   56969 => x"7C",
						   -- Begin: __mspabi_slli_12
						   56970 => x"0C",		-- 00de8a: 0C5C             RLA.W   R12
						   56971 => x"7C",
						   -- Begin: __mspabi_slli_11
						   56972 => x"0C",		-- 00de8c: 0C5C             RLA.W   R12
						   56973 => x"7C",
						   -- Begin: __mspabi_slli_10
						   56974 => x"0C",		-- 00de8e: 0C5C             RLA.W   R12
						   56975 => x"7C",
						   -- Begin: __mspabi_slli_9
						   56976 => x"0C",		-- 00de90: 0C5C             RLA.W   R12
						   56977 => x"7C",
						   -- Begin: __mspabi_slli_8
						   56978 => x"0C",		-- 00de92: 0C5C             RLA.W   R12
						   56979 => x"7C",
						   -- Begin: __mspabi_slli_7
						   56980 => x"0C",		-- 00de94: 0C5C             RLA.W   R12
						   56981 => x"7C",
						   -- Begin: __mspabi_slli_6
						   56982 => x"0C",		-- 00de96: 0C5C             RLA.W   R12
						   56983 => x"7C",
						   -- Begin: __mspabi_slli_5
						   56984 => x"0C",		-- 00de98: 0C5C             RLA.W   R12
						   56985 => x"7C",
						   -- Begin: __mspabi_slli_4
						   56986 => x"0C",		-- 00de9a: 0C5C             RLA.W   R12
						   56987 => x"7C",
						   -- Begin: __mspabi_slli_3
						   56988 => x"0C",		-- 00de9c: 0C5C             RLA.W   R12
						   56989 => x"7C",
						   -- Begin: __mspabi_slli_2
						   56990 => x"0C",		-- 00de9e: 0C5C             RLA.W   R12
						   56991 => x"7C",
						   -- Begin: __mspabi_slli_1
						   56992 => x"0C",		-- 00dea0: 0C5C             RLA.W   R12
						   56993 => x"7C",
						   56994 => x"30",		-- 00dea2: 3041             RET     
						   56995 => x"61",
						   -- Begin: strncpy
						   56996 => x"0E",		-- 00dea4: 0E93             TST.W   R14
						   56997 => x"B3",
						   56998 => x"13",		-- 00dea6: 1324             JEQ     ($C$L4)
						   56999 => x"44",
						   57000 => x"0F",		-- 00dea8: 0F4C             MOV.W   R12,R15
						   57001 => x"6C",
						   57002 => x"6B",		-- 00deaa: 6B4D             MOV.B   @R13,R11
						   57003 => x"6D",
						   57004 => x"1F",		-- 00deac: 1F53             INC.W   R15
						   57005 => x"73",
						   57006 => x"CF",		-- 00deae: CF4B             MOV.B   R11,0xffff(R15)
						   57007 => x"6B",
						   57008 => x"FF",		-- 00deb0: FFFF            
						   57009 => x"FF",
						   57010 => x"0B",		-- 00deb2: 0B93             TST.W   R11
						   57011 => x"B3",
						   57012 => x"03",		-- 00deb4: 0324             JEQ     ($C$L2)
						   57013 => x"44",
						   57014 => x"1D",		-- 00deb6: 1D53             INC.W   R13
						   57015 => x"73",
						   57016 => x"1E",		-- 00deb8: 1E83             DEC.W   R14
						   57017 => x"A3",
						   57018 => x"F7",		-- 00deba: F723             JNE     ($C$L1)
						   57019 => x"43",
						   57020 => x"0D",		-- 00debc: 0D4E             MOV.W   R14,R13
						   57021 => x"6E",
						   57022 => x"1E",		-- 00debe: 1E83             DEC.W   R14
						   57023 => x"A3",
						   57024 => x"2D",		-- 00dec0: 2D93             CMP.W   #2,R13
						   57025 => x"B3",
						   57026 => x"05",		-- 00dec2: 0528             JLO     ($C$L4)
						   57027 => x"48",
						   57028 => x"1F",		-- 00dec4: 1F53             INC.W   R15
						   57029 => x"73",
						   57030 => x"CF",		-- 00dec6: CF43             CLR.B   0xffff(R15)
						   57031 => x"63",
						   57032 => x"FF",		-- 00dec8: FFFF            
						   57033 => x"FF",
						   57034 => x"1E",		-- 00deca: 1E83             DEC.W   R14
						   57035 => x"A3",
						   57036 => x"FB",		-- 00decc: FB23             JNE     ($C$L3)
						   57037 => x"43",
						   57038 => x"30",		-- 00dece: 3041             RET     
						   57039 => x"61",
						   -- Begin: __mspabi_negd
						   57040 => x"31",		-- 00ded0: 3182             SUB.W   #8,SP
						   57041 => x"A2",
						   57042 => x"81",		-- 00ded2: 814C             MOV.W   R12,0x0000(SP)
						   57043 => x"6C",
						   57044 => x"00",		-- 00ded4: 0000            
						   57045 => x"00",
						   57046 => x"81",		-- 00ded6: 814D             MOV.W   R13,0x0002(SP)
						   57047 => x"6D",
						   57048 => x"02",		-- 00ded8: 0200            
						   57049 => x"00",
						   57050 => x"81",		-- 00deda: 814E             MOV.W   R14,0x0004(SP)
						   57051 => x"6E",
						   57052 => x"04",		-- 00dedc: 0400            
						   57053 => x"00",
						   57054 => x"81",		-- 00dede: 814F             MOV.W   R15,0x0006(SP)
						   57055 => x"6F",
						   57056 => x"06",		-- 00dee0: 0600            
						   57057 => x"00",
						   57058 => x"F1",		-- 00dee2: F1E0             XOR.B   #0x0080,0x0007(SP)
						   57059 => x"00",
						   57060 => x"80",		-- 00dee4: 8000            
						   57061 => x"00",
						   57062 => x"07",		-- 00dee6: 0700            
						   57063 => x"00",
						   57064 => x"2C",		-- 00dee8: 2C41             MOV.W   @SP,R12
						   57065 => x"61",
						   57066 => x"1D",		-- 00deea: 1D41             MOV.W   0x0002(SP),R13
						   57067 => x"61",
						   57068 => x"02",		-- 00deec: 0200            
						   57069 => x"00",
						   57070 => x"1E",		-- 00deee: 1E41             MOV.W   0x0004(SP),R14
						   57071 => x"61",
						   57072 => x"04",		-- 00def0: 0400            
						   57073 => x"00",
						   57074 => x"1F",		-- 00def2: 1F41             MOV.W   0x0006(SP),R15
						   57075 => x"61",
						   57076 => x"06",		-- 00def4: 0600            
						   57077 => x"00",
						   57078 => x"31",		-- 00def6: 3152             ADD.W   #8,SP
						   57079 => x"72",
						   57080 => x"30",		-- 00def8: 3041             RET     
						   57081 => x"61",
						   -- Begin: __mspabi_fixdi
						   57082 => x"B0",		-- 00defa: B012             CALL    #__mspabi_fixdli
						   57083 => x"32",
						   57084 => x"9A",		-- 00defc: 9AD4            
						   57085 => x"D4",
						   57086 => x"0D",		-- 00defe: 0D93             TST.W   R13
						   57087 => x"B3",
						   57088 => x"07",		-- 00df00: 0738             JL      ($C$L7)
						   57089 => x"58",
						   57090 => x"03",		-- 00df02: 0320             JNE     ($C$L6)
						   57091 => x"40",
						   57092 => x"3C",		-- 00df04: 3C90             CMP.W   #0x8000,R12
						   57093 => x"B0",
						   57094 => x"00",		-- 00df06: 0080            
						   57095 => x"80",
						   57096 => x"03",		-- 00df08: 0328             JLO     ($C$L7)
						   57097 => x"48",
						   57098 => x"3C",		-- 00df0a: 3C40             MOV.W   #0x7fff,R12
						   57099 => x"60",
						   57100 => x"FF",		-- 00df0c: FF7F            
						   57101 => x"7F",
						   57102 => x"30",		-- 00df0e: 3041             RET     
						   57103 => x"61",
						   57104 => x"3D",		-- 00df10: 3D93             CMP.W   #-1,R13
						   57105 => x"B3",
						   57106 => x"04",		-- 00df12: 0438             JL      ($C$L8)
						   57107 => x"58",
						   57108 => x"05",		-- 00df14: 0520             JNE     ($C$L9)
						   57109 => x"40",
						   57110 => x"3C",		-- 00df16: 3C90             CMP.W   #0x8000,R12
						   57111 => x"B0",
						   57112 => x"00",		-- 00df18: 0080            
						   57113 => x"80",
						   57114 => x"02",		-- 00df1a: 022C             JHS     ($C$L9)
						   57115 => x"4C",
						   57116 => x"3C",		-- 00df1c: 3C40             MOV.W   #0x8000,R12
						   57117 => x"60",
						   57118 => x"00",		-- 00df1e: 0080            
						   57119 => x"80",
						   57120 => x"30",		-- 00df20: 3041             RET     
						   57121 => x"61",
						   -- Begin: free_list_insert
						   57122 => x"2F",		-- 00df22: 2F4C             MOV.W   @R12,R15
						   57123 => x"6C",
						   57124 => x"1F",		-- 00df24: 1FC3             BIC.W   #1,R15
						   57125 => x"E3",
						   57126 => x"3E",		-- 00df26: 3E40             MOV.W   #0x21a6,R14
						   57127 => x"60",
						   57128 => x"A6",		-- 00df28: A621            
						   57129 => x"21",
						   57130 => x"03",		-- 00df2a: 033C             JMP     ($C$L5)
						   57131 => x"5C",
						   57132 => x"2D",		-- 00df2c: 2D42             MOV.W   #4,R13
						   57133 => x"62",
						   57134 => x"2D",		-- 00df2e: 2D5E             ADD.W   @R14,R13
						   57135 => x"7E",
						   57136 => x"0E",		-- 00df30: 0E4D             MOV.W   R13,R14
						   57137 => x"6D",
						   57138 => x"2D",		-- 00df32: 2D4E             MOV.W   @R14,R13
						   57139 => x"6E",
						   57140 => x"0D",		-- 00df34: 0D93             TST.W   R13
						   57141 => x"B3",
						   57142 => x"04",		-- 00df36: 0424             JEQ     ($C$L6)
						   57143 => x"44",
						   57144 => x"2D",		-- 00df38: 2D4D             MOV.W   @R13,R13
						   57145 => x"6D",
						   57146 => x"1D",		-- 00df3a: 1DC3             BIC.W   #1,R13
						   57147 => x"E3",
						   57148 => x"0D",		-- 00df3c: 0D9F             CMP.W   R15,R13
						   57149 => x"BF",
						   57150 => x"F6",		-- 00df3e: F62B             JLO     ($C$L4)
						   57151 => x"4B",
						   57152 => x"AC",		-- 00df40: AC4E             MOV.W   @R14,0x0004(R12)
						   57153 => x"6E",
						   57154 => x"04",		-- 00df42: 0400            
						   57155 => x"00",
						   57156 => x"8E",		-- 00df44: 8E4C             MOV.W   R12,0x0000(R14)
						   57157 => x"6C",
						   57158 => x"00",		-- 00df46: 0000            
						   57159 => x"00",
						   57160 => x"30",		-- 00df48: 3041             RET     
						   57161 => x"61",
						   -- Begin: remove
						   -- Begin: unlink
						   57162 => x"0A",		-- 00df4a: 0A12             PUSH    R10
						   57163 => x"32",
						   57164 => x"21",		-- 00df4c: 2183             DECD.W  SP
						   57165 => x"A3",
						   57166 => x"81",		-- 00df4e: 814C             MOV.W   R12,0x0000(SP)
						   57167 => x"6C",
						   57168 => x"00",		-- 00df50: 0000            
						   57169 => x"00",
						   57170 => x"92",		-- 00df52: 9212             CALL    &_lock
						   57171 => x"32",
						   57172 => x"F2",		-- 00df54: F220            
						   57173 => x"20",
						   57174 => x"0C",		-- 00df56: 0C41             MOV.W   SP,R12
						   57175 => x"61",
						   57176 => x"B0",		-- 00df58: B012             CALL    #getdevice
						   57177 => x"32",
						   57178 => x"34",		-- 00df5a: 34D8            
						   57179 => x"D8",
						   57180 => x"0F",		-- 00df5c: 0F4C             MOV.W   R12,R15
						   57181 => x"6C",
						   57182 => x"2C",		-- 00df5e: 2C41             MOV.W   @SP,R12
						   57183 => x"61",
						   57184 => x"9F",		-- 00df60: 9F12             CALL    0x0016(R15)
						   57185 => x"32",
						   57186 => x"16",		-- 00df62: 1600            
						   57187 => x"00",
						   57188 => x"0A",		-- 00df64: 0A4C             MOV.W   R12,R10
						   57189 => x"6C",
						   57190 => x"92",		-- 00df66: 9212             CALL    &_unlock
						   57191 => x"32",
						   57192 => x"F4",		-- 00df68: F420            
						   57193 => x"20",
						   57194 => x"0C",		-- 00df6a: 0C4A             MOV.W   R10,R12
						   57195 => x"6A",
						   57196 => x"21",		-- 00df6c: 2153             INCD.W  SP
						   57197 => x"73",
						   57198 => x"3A",		-- 00df6e: 3A41             POP.W   R10
						   57199 => x"61",
						   57200 => x"30",		-- 00df70: 3041             RET     
						   57201 => x"61",
						   -- Begin: lseek
						   57202 => x"0C",		-- 00df72: 0C93             TST.W   R12
						   57203 => x"B3",
						   57204 => x"0E",		-- 00df74: 0E38             JL      ($C$L1)
						   57205 => x"58",
						   57206 => x"3C",		-- 00df76: 3C90             CMP.W   #0x000a,R12
						   57207 => x"B0",
						   57208 => x"0A",		-- 00df78: 0A00            
						   57209 => x"00",
						   57210 => x"0B",		-- 00df7a: 0B34             JGE     ($C$L1)
						   57211 => x"54",
						   57212 => x"0C",		-- 00df7c: 0C5C             RLA.W   R12
						   57213 => x"7C",
						   57214 => x"0C",		-- 00df7e: 0C5C             RLA.W   R12
						   57215 => x"7C",
						   57216 => x"3C",		-- 00df80: 3C50             ADD.W   #0x20c6,R12
						   57217 => x"70",
						   57218 => x"C6",		-- 00df82: C620            
						   57219 => x"20",
						   57220 => x"2B",		-- 00df84: 2B4C             MOV.W   @R12,R11
						   57221 => x"6C",
						   57222 => x"0B",		-- 00df86: 0B93             TST.W   R11
						   57223 => x"B3",
						   57224 => x"04",		-- 00df88: 0424             JEQ     ($C$L1)
						   57225 => x"44",
						   57226 => x"1C",		-- 00df8a: 1C4C             MOV.W   0x0002(R12),R12
						   57227 => x"6C",
						   57228 => x"02",		-- 00df8c: 0200            
						   57229 => x"00",
						   57230 => x"10",		-- 00df8e: 104B             BR      0x0014(R11)
						   57231 => x"6B",
						   57232 => x"14",		-- 00df90: 1400            
						   57233 => x"00",
						   57234 => x"3C",		-- 00df92: 3C43             MOV.W   #-1,R12
						   57235 => x"63",
						   57236 => x"3D",		-- 00df94: 3D43             MOV.W   #-1,R13
						   57237 => x"63",
						   57238 => x"30",		-- 00df96: 3041             RET     
						   57239 => x"61",
						   -- Begin: __mspabi_mpyl
						   -- Begin: __mspabi_mpyl_sw
						   57240 => x"0A",		-- 00df98: 0A12             PUSH    R10
						   57241 => x"32",
						   57242 => x"0A",		-- 00df9a: 0A43             CLR.W   R10
						   57243 => x"63",
						   57244 => x"0B",		-- 00df9c: 0B43             CLR.W   R11
						   57245 => x"63",
						   -- Begin: mpyl_add_loop
						   57246 => x"12",		-- 00df9e: 12C3             CLRC    
						   57247 => x"E3",
						   57248 => x"0D",		-- 00dfa0: 0D10             RRC     R13
						   57249 => x"30",
						   57250 => x"0C",		-- 00dfa2: 0C10             RRC     R12
						   57251 => x"30",
						   57252 => x"02",		-- 00dfa4: 0228             JLO     (shift_test_mpyl)
						   57253 => x"48",
						   57254 => x"0A",		-- 00dfa6: 0A5E             ADD.W   R14,R10
						   57255 => x"7E",
						   57256 => x"0B",		-- 00dfa8: 0B6F             ADDC.W  R15,R11
						   57257 => x"8F",
						   -- Begin: shift_test_mpyl
						   57258 => x"0E",		-- 00dfaa: 0E5E             RLA.W   R14
						   57259 => x"7E",
						   57260 => x"0F",		-- 00dfac: 0F6F             RLC.W   R15
						   57261 => x"8F",
						   57262 => x"0D",		-- 00dfae: 0D93             TST.W   R13
						   57263 => x"B3",
						   57264 => x"F6",		-- 00dfb0: F623             JNE     (mpyl_add_loop)
						   57265 => x"43",
						   57266 => x"0C",		-- 00dfb2: 0C93             TST.W   R12
						   57267 => x"B3",
						   57268 => x"F4",		-- 00dfb4: F423             JNE     (mpyl_add_loop)
						   57269 => x"43",
						   57270 => x"0C",		-- 00dfb6: 0C4A             MOV.W   R10,R12
						   57271 => x"6A",
						   57272 => x"0D",		-- 00dfb8: 0D4B             MOV.W   R11,R13
						   57273 => x"6B",
						   57274 => x"3A",		-- 00dfba: 3A41             POP.W   R10
						   57275 => x"61",
						   57276 => x"30",		-- 00dfbc: 3041             RET     
						   57277 => x"61",
						   -- Begin: write
						   57278 => x"0C",		-- 00dfbe: 0C93             TST.W   R12
						   57279 => x"B3",
						   57280 => x"0E",		-- 00dfc0: 0E38             JL      ($C$L1)
						   57281 => x"58",
						   57282 => x"3C",		-- 00dfc2: 3C90             CMP.W   #0x000a,R12
						   57283 => x"B0",
						   57284 => x"0A",		-- 00dfc4: 0A00            
						   57285 => x"00",
						   57286 => x"0B",		-- 00dfc6: 0B34             JGE     ($C$L1)
						   57287 => x"54",
						   57288 => x"0C",		-- 00dfc8: 0C5C             RLA.W   R12
						   57289 => x"7C",
						   57290 => x"0C",		-- 00dfca: 0C5C             RLA.W   R12
						   57291 => x"7C",
						   57292 => x"3C",		-- 00dfcc: 3C50             ADD.W   #0x20c6,R12
						   57293 => x"70",
						   57294 => x"C6",		-- 00dfce: C620            
						   57295 => x"20",
						   57296 => x"2F",		-- 00dfd0: 2F4C             MOV.W   @R12,R15
						   57297 => x"6C",
						   57298 => x"0F",		-- 00dfd2: 0F93             TST.W   R15
						   57299 => x"B3",
						   57300 => x"04",		-- 00dfd4: 0424             JEQ     ($C$L1)
						   57301 => x"44",
						   57302 => x"1C",		-- 00dfd6: 1C4C             MOV.W   0x0002(R12),R12
						   57303 => x"6C",
						   57304 => x"02",		-- 00dfd8: 0200            
						   57305 => x"00",
						   57306 => x"10",		-- 00dfda: 104F             BR      0x0012(R15)
						   57307 => x"6F",
						   57308 => x"12",		-- 00dfdc: 1200            
						   57309 => x"00",
						   57310 => x"3C",		-- 00dfde: 3C43             MOV.W   #-1,R12
						   57311 => x"63",
						   57312 => x"30",		-- 00dfe0: 3041             RET     
						   57313 => x"61",
						   -- Begin: __mspabi_mpyul
						   -- Begin: __mspabi_mpyul_sw
						   57314 => x"0B",		-- 00dfe2: 0B4C             MOV.W   R12,R11
						   57315 => x"6C",
						   57316 => x"0E",		-- 00dfe4: 0E4D             MOV.W   R13,R14
						   57317 => x"6D",
						   57318 => x"0F",		-- 00dfe6: 0F43             CLR.W   R15
						   57319 => x"63",
						   57320 => x"0C",		-- 00dfe8: 0C43             CLR.W   R12
						   57321 => x"63",
						   57322 => x"0D",		-- 00dfea: 0D43             CLR.W   R13
						   57323 => x"63",
						   57324 => x"12",		-- 00dfec: 12C3             CLRC    
						   57325 => x"E3",
						   57326 => x"0B",		-- 00dfee: 0B10             RRC     R11
						   57327 => x"30",
						   57328 => x"01",		-- 00dff0: 013C             JMP     (mpyul_add_loop1)
						   57329 => x"5C",
						   -- Begin: mpyul_add_loop
						   57330 => x"0B",		-- 00dff2: 0B11             RRA     R11
						   57331 => x"31",
						   -- Begin: mpyul_add_loop1
						   57332 => x"02",		-- 00dff4: 0228             JLO     (shift_test_mpyul)
						   57333 => x"48",
						   57334 => x"0C",		-- 00dff6: 0C5E             ADD.W   R14,R12
						   57335 => x"7E",
						   57336 => x"0D",		-- 00dff8: 0D6F             ADDC.W  R15,R13
						   57337 => x"8F",
						   -- Begin: shift_test_mpyul
						   57338 => x"0E",		-- 00dffa: 0E5E             RLA.W   R14
						   57339 => x"7E",
						   57340 => x"0F",		-- 00dffc: 0F6F             RLC.W   R15
						   57341 => x"8F",
						   57342 => x"0B",		-- 00dffe: 0B93             TST.W   R11
						   57343 => x"B3",
						   57344 => x"F8",		-- 00e000: F823             JNE     (mpyul_add_loop)
						   57345 => x"43",
						   57346 => x"30",		-- 00e002: 3041             RET     
						   57347 => x"61",
						   -- Begin: memccpy
						   57348 => x"0A",		-- 00e004: 0A12             PUSH    R10
						   57349 => x"32",
						   57350 => x"0F",		-- 00e006: 0F93             TST.W   R15
						   57351 => x"B3",
						   57352 => x"0B",		-- 00e008: 0B24             JEQ     ($C$L2)
						   57353 => x"44",
						   57354 => x"4E",		-- 00e00a: 4E4E             MOV.B   R14,R14
						   57355 => x"6E",
						   57356 => x"6B",		-- 00e00c: 6B4D             MOV.B   @R13,R11
						   57357 => x"6D",
						   57358 => x"1C",		-- 00e00e: 1C53             INC.W   R12
						   57359 => x"73",
						   57360 => x"CC",		-- 00e010: CC4B             MOV.B   R11,0xffff(R12)
						   57361 => x"6B",
						   57362 => x"FF",		-- 00e012: FFFF            
						   57363 => x"FF",
						   57364 => x"4A",		-- 00e014: 4A4E             MOV.B   R14,R10
						   57365 => x"6E",
						   57366 => x"0B",		-- 00e016: 0B9A             CMP.W   R10,R11
						   57367 => x"BA",
						   57368 => x"04",		-- 00e018: 0424             JEQ     ($C$L3)
						   57369 => x"44",
						   57370 => x"1D",		-- 00e01a: 1D53             INC.W   R13
						   57371 => x"73",
						   57372 => x"1F",		-- 00e01c: 1F83             DEC.W   R15
						   57373 => x"A3",
						   57374 => x"F6",		-- 00e01e: F623             JNE     ($C$L1)
						   57375 => x"43",
						   57376 => x"0C",		-- 00e020: 0C43             CLR.W   R12
						   57377 => x"63",
						   57378 => x"3A",		-- 00e022: 3A41             POP.W   R10
						   57379 => x"61",
						   57380 => x"30",		-- 00e024: 3041             RET     
						   57381 => x"61",
						   -- Begin: __mspabi_mpyull
						   -- Begin: __mspabi_mpyull_sw
						   57382 => x"0A",		-- 00e026: 0A12             PUSH    R10
						   57383 => x"32",
						   57384 => x"09",		-- 00e028: 0912             PUSH    R9
						   57385 => x"32",
						   57386 => x"08",		-- 00e02a: 0812             PUSH    R8
						   57387 => x"32",
						   57388 => x"08",		-- 00e02c: 084C             MOV.W   R12,R8
						   57389 => x"6C",
						   57390 => x"09",		-- 00e02e: 094D             MOV.W   R13,R9
						   57391 => x"6D",
						   57392 => x"0A",		-- 00e030: 0A43             CLR.W   R10
						   57393 => x"63",
						   57394 => x"0B",		-- 00e032: 0B43             CLR.W   R11
						   57395 => x"63",
						   57396 => x"0C",		-- 00e034: 0C4E             MOV.W   R14,R12
						   57397 => x"6E",
						   57398 => x"0D",		-- 00e036: 0D4F             MOV.W   R15,R13
						   57399 => x"6F",
						   57400 => x"0E",		-- 00e038: 0E43             CLR.W   R14
						   57401 => x"63",
						   57402 => x"0F",		-- 00e03a: 0F43             CLR.W   R15
						   57403 => x"63",
						   57404 => x"B0",		-- 00e03c: B012             CALL    #__mspabi_mpyll_sw
						   57405 => x"32",
						   57406 => x"E6",		-- 00e03e: E6C5            
						   57407 => x"C5",
						   57408 => x"30",		-- 00e040: 3040             BR      #__mspabi_func_epilog_3
						   57409 => x"60",
						   57410 => x"78",		-- 00e042: 78E1            
						   57411 => x"E1",
						   -- Begin: _c_int00_noargs
						   57412 => x"31",		-- 00e044: 3140             MOV.W   #0x3000,SP
						   57413 => x"60",
						   57414 => x"00",		-- 00e046: 0030            
						   57415 => x"30",
						   57416 => x"B0",		-- 00e048: B012             CALL    #_system_pre_init
						   57417 => x"32",
						   57418 => x"D8",		-- 00e04a: D8E1            
						   57419 => x"E1",
						   57420 => x"0C",		-- 00e04c: 0C93             TST.W   R12
						   57421 => x"B3",
						   57422 => x"02",		-- 00e04e: 0224             JEQ     ($C$L2)
						   57423 => x"44",
						   57424 => x"B0",		-- 00e050: B012             CALL    #__TI_auto_init_nobinit_nopinit
						   57425 => x"32",
						   57426 => x"76",		-- 00e052: 76DB            
						   57427 => x"DB",
						   57428 => x"0C",		-- 00e054: 0C43             CLR.W   R12
						   57429 => x"63",
						   57430 => x"B0",		-- 00e056: B012             CALL    #main
						   57431 => x"32",
						   57432 => x"B4",		-- 00e058: B4DC            
						   57433 => x"DC",
						   57434 => x"1C",		-- 00e05a: 1C43             MOV.W   #1,R12
						   57435 => x"63",
						   57436 => x"B0",		-- 00e05c: B012             CALL    #exit
						   57437 => x"32",
						   57438 => x"32",		-- 00e05e: 32DB            
						   57439 => x"DB",
						   -- Begin: free_list_remove
						   57440 => x"3F",		-- 00e060: 3F40             MOV.W   #0x21a6,R15
						   57441 => x"60",
						   57442 => x"A6",		-- 00e062: A621            
						   57443 => x"21",
						   57444 => x"02",		-- 00e064: 023C             JMP     ($C$L2)
						   57445 => x"5C",
						   57446 => x"2F",		-- 00e066: 2F42             MOV.W   #4,R15
						   57447 => x"62",
						   57448 => x"0F",		-- 00e068: 0F5E             ADD.W   R14,R15
						   57449 => x"7E",
						   57450 => x"2E",		-- 00e06a: 2E4F             MOV.W   @R15,R14
						   57451 => x"6F",
						   57452 => x"0E",		-- 00e06c: 0E93             TST.W   R14
						   57453 => x"B3",
						   57454 => x"05",		-- 00e06e: 0524             JEQ     ($C$L3)
						   57455 => x"44",
						   57456 => x"0E",		-- 00e070: 0E9C             CMP.W   R12,R14
						   57457 => x"BC",
						   57458 => x"F9",		-- 00e072: F923             JNE     ($C$L1)
						   57459 => x"43",
						   57460 => x"9F",		-- 00e074: 9F4C             MOV.W   0x0004(R12),0x0000(R15)
						   57461 => x"6C",
						   57462 => x"04",		-- 00e076: 0400            
						   57463 => x"00",
						   57464 => x"00",		-- 00e078: 0000            
						   57465 => x"00",
						   57466 => x"30",		-- 00e07a: 3041             RET     
						   57467 => x"61",
						   -- Begin: strchr
						   57468 => x"6F",		-- 00e07c: 6F4C             MOV.B   @R12,R15
						   57469 => x"6C",
						   57470 => x"4D",		-- 00e07e: 4D4D             MOV.B   R13,R13
						   57471 => x"6D",
						   57472 => x"06",		-- 00e080: 063C             JMP     ($C$L3)
						   57473 => x"5C",
						   57474 => x"0F",		-- 00e082: 0F93             TST.W   R15
						   57475 => x"B3",
						   57476 => x"02",		-- 00e084: 0220             JNE     ($C$L2)
						   57477 => x"40",
						   57478 => x"0C",		-- 00e086: 0C43             CLR.W   R12
						   57479 => x"63",
						   57480 => x"30",		-- 00e088: 3041             RET     
						   57481 => x"61",
						   57482 => x"1C",		-- 00e08a: 1C53             INC.W   R12
						   57483 => x"73",
						   57484 => x"6F",		-- 00e08c: 6F4C             MOV.B   @R12,R15
						   57485 => x"6C",
						   57486 => x"4E",		-- 00e08e: 4E4D             MOV.B   R13,R14
						   57487 => x"6D",
						   57488 => x"0F",		-- 00e090: 0F9E             CMP.W   R14,R15
						   57489 => x"BE",
						   57490 => x"F7",		-- 00e092: F723             JNE     ($C$L1)
						   57491 => x"43",
						   57492 => x"30",		-- 00e094: 3041             RET     
						   57493 => x"61",
						   -- Begin: strcmp
						   57494 => x"0F",		-- 00e096: 0F4C             MOV.W   R12,R15
						   57495 => x"6C",
						   57496 => x"6E",		-- 00e098: 6E4F             MOV.B   @R15,R14
						   57497 => x"6F",
						   57498 => x"6B",		-- 00e09a: 6B4D             MOV.B   @R13,R11
						   57499 => x"6D",
						   57500 => x"4C",		-- 00e09c: 4C4E             MOV.B   R14,R12
						   57501 => x"6E",
						   57502 => x"0C",		-- 00e09e: 0C8B             SUB.W   R11,R12
						   57503 => x"AB",
						   57504 => x"4E",		-- 00e0a0: 4E93             TST.B   R14
						   57505 => x"B3",
						   57506 => x"04",		-- 00e0a2: 0424             JEQ     ($C$L2)
						   57507 => x"44",
						   57508 => x"1D",		-- 00e0a4: 1D53             INC.W   R13
						   57509 => x"73",
						   57510 => x"1F",		-- 00e0a6: 1F53             INC.W   R15
						   57511 => x"73",
						   57512 => x"0C",		-- 00e0a8: 0C93             TST.W   R12
						   57513 => x"B3",
						   57514 => x"F6",		-- 00e0aa: F627             JEQ     ($C$L1)
						   57515 => x"47",
						   57516 => x"30",		-- 00e0ac: 3041             RET     
						   57517 => x"61",
						   -- Begin: __mspabi_divu
						   -- Begin: __mspabi_remu
						   57518 => x"0E",		-- 00e0ae: 0E43             CLR.W   R14
						   57519 => x"63",
						   57520 => x"0F",		-- 00e0b0: 0F4C             MOV.W   R12,R15
						   57521 => x"6C",
						   57522 => x"1C",		-- 00e0b2: 1C43             MOV.W   #1,R12
						   57523 => x"63",
						   -- Begin: div_loop
						   57524 => x"0F",		-- 00e0b4: 0F5F             RLA.W   R15
						   57525 => x"7F",
						   57526 => x"0E",		-- 00e0b6: 0E6E             RLC.W   R14
						   57527 => x"8E",
						   57528 => x"0E",		-- 00e0b8: 0E9D             CMP.W   R13,R14
						   57529 => x"BD",
						   57530 => x"01",		-- 00e0ba: 0128             JLO     (set_quotient_bit)
						   57531 => x"48",
						   57532 => x"0E",		-- 00e0bc: 0E8D             SUB.W   R13,R14
						   57533 => x"AD",
						   -- Begin: set_quotient_bit
						   57534 => x"0C",		-- 00e0be: 0C6C             RLC.W   R12
						   57535 => x"8C",
						   57536 => x"F9",		-- 00e0c0: F92B             JLO     (div_loop)
						   57537 => x"4B",
						   57538 => x"30",		-- 00e0c2: 3041             RET     
						   57539 => x"61",
						   -- Begin: __TI_zero_init_nomemset
						   57540 => x"1F",		-- 00e0c4: 1F4C             MOV.W   0x0001(R12),R15
						   57541 => x"6C",
						   57542 => x"01",		-- 00e0c6: 0100            
						   57543 => x"00",
						   57544 => x"0F",		-- 00e0c8: 0F93             TST.W   R15
						   57545 => x"B3",
						   57546 => x"05",		-- 00e0ca: 0524             JEQ     ($C$L2)
						   57547 => x"44",
						   57548 => x"1D",		-- 00e0cc: 1D53             INC.W   R13
						   57549 => x"73",
						   57550 => x"CD",		-- 00e0ce: CD43             CLR.B   0xffff(R13)
						   57551 => x"63",
						   57552 => x"FF",		-- 00e0d0: FFFF            
						   57553 => x"FF",
						   57554 => x"1F",		-- 00e0d2: 1F83             DEC.W   R15
						   57555 => x"A3",
						   57556 => x"FB",		-- 00e0d4: FB23             JNE     ($C$L1)
						   57557 => x"43",
						   57558 => x"30",		-- 00e0d6: 3041             RET     
						   57559 => x"61",
						   -- Begin: memchr
						   57560 => x"0E",		-- 00e0d8: 0E93             TST.W   R14
						   57561 => x"B3",
						   57562 => x"06",		-- 00e0da: 0624             JEQ     ($C$L2)
						   57563 => x"44",
						   57564 => x"4D",		-- 00e0dc: 4D4D             MOV.B   R13,R13
						   57565 => x"6D",
						   57566 => x"6D",		-- 00e0de: 6D9C             CMP.B   @R12,R13
						   57567 => x"BC",
						   57568 => x"04",		-- 00e0e0: 0424             JEQ     ($C$L3)
						   57569 => x"44",
						   57570 => x"1C",		-- 00e0e2: 1C53             INC.W   R12
						   57571 => x"73",
						   57572 => x"1E",		-- 00e0e4: 1E83             DEC.W   R14
						   57573 => x"A3",
						   57574 => x"FB",		-- 00e0e6: FB23             JNE     ($C$L1)
						   57575 => x"43",
						   57576 => x"0C",		-- 00e0e8: 0C43             CLR.W   R12
						   57577 => x"63",
						   57578 => x"30",		-- 00e0ea: 3041             RET     
						   57579 => x"61",
						   -- Begin: memset
						   57580 => x"0F",		-- 00e0ec: 0F4C             MOV.W   R12,R15
						   57581 => x"6C",
						   57582 => x"0E",		-- 00e0ee: 0E93             TST.W   R14
						   57583 => x"B3",
						   57584 => x"06",		-- 00e0f0: 0624             JEQ     ($C$L2)
						   57585 => x"44",
						   57586 => x"4D",		-- 00e0f2: 4D4D             MOV.B   R13,R13
						   57587 => x"6D",
						   57588 => x"1F",		-- 00e0f4: 1F53             INC.W   R15
						   57589 => x"73",
						   57590 => x"CF",		-- 00e0f6: CF4D             MOV.B   R13,0xffff(R15)
						   57591 => x"6D",
						   57592 => x"FF",		-- 00e0f8: FFFF            
						   57593 => x"FF",
						   57594 => x"1E",		-- 00e0fa: 1E83             DEC.W   R14
						   57595 => x"A3",
						   57596 => x"FB",		-- 00e0fc: FB23             JNE     ($C$L1)
						   57597 => x"43",
						   57598 => x"30",		-- 00e0fe: 3041             RET     
						   57599 => x"61",
						   -- Begin: __mspabi_mpyi
						   -- Begin: __mspabi_mpyi_sw
						   57600 => x"0E",		-- 00e100: 0E43             CLR.W   R14
						   57601 => x"63",
						   -- Begin: mpyi_add_loop
						   57602 => x"12",		-- 00e102: 12C3             CLRC    
						   57603 => x"E3",
						   57604 => x"0C",		-- 00e104: 0C10             RRC     R12
						   57605 => x"30",
						   57606 => x"01",		-- 00e106: 0128             JLO     (shift_test_mpyi)
						   57607 => x"48",
						   57608 => x"0E",		-- 00e108: 0E5D             ADD.W   R13,R14
						   57609 => x"7D",
						   -- Begin: shift_test_mpyi
						   57610 => x"0D",		-- 00e10a: 0D5D             RLA.W   R13
						   57611 => x"7D",
						   57612 => x"0C",		-- 00e10c: 0C93             TST.W   R12
						   57613 => x"B3",
						   57614 => x"F9",		-- 00e10e: F923             JNE     (mpyi_add_loop)
						   57615 => x"43",
						   57616 => x"0C",		-- 00e110: 0C4E             MOV.W   R14,R12
						   57617 => x"6E",
						   57618 => x"30",		-- 00e112: 3041             RET     
						   57619 => x"61",
						   -- Begin: wcslen
						   57620 => x"0F",		-- 00e114: 0F4C             MOV.W   R12,R15
						   57621 => x"6C",
						   57622 => x"01",		-- 00e116: 013C             JMP     ($C$L2)
						   57623 => x"5C",
						   57624 => x"2F",		-- 00e118: 2F53             INCD.W  R15
						   57625 => x"73",
						   57626 => x"8F",		-- 00e11a: 8F93             TST.W   0x0000(R15)
						   57627 => x"B3",
						   57628 => x"00",		-- 00e11c: 0000            
						   57629 => x"00",
						   57630 => x"FC",		-- 00e11e: FC23             JNE     ($C$L1)
						   57631 => x"43",
						   57632 => x"0F",		-- 00e120: 0F8C             SUB.W   R12,R15
						   57633 => x"AC",
						   57634 => x"0F",		-- 00e122: 0F11             RRA     R15
						   57635 => x"31",
						   57636 => x"0C",		-- 00e124: 0C4F             MOV.W   R15,R12
						   57637 => x"6F",
						   57638 => x"30",		-- 00e126: 3041             RET     
						   57639 => x"61",
						   -- Begin: buff_value
						   57640 => x"21",		-- 00e128: 2183             DECD.W  SP
						   57641 => x"A3",
						   57642 => x"81",		-- 00e12a: 814C             MOV.W   R12,0x0000(SP)
						   57643 => x"6C",
						   57644 => x"00",		-- 00e12c: 0000            
						   57645 => x"00",
						   57646 => x"3D",		-- 00e12e: 3D40             MOV.W   #0x8514,R13
						   57647 => x"60",
						   57648 => x"14",		-- 00e130: 1485            
						   57649 => x"85",
						   57650 => x"B0",		-- 00e132: B012             CALL    #strcpy
						   57651 => x"32",
						   57652 => x"80",		-- 00e134: 80E1            
						   57653 => x"E1",
						   57654 => x"21",		-- 00e136: 2153             INCD.W  SP
						   57655 => x"73",
						   57656 => x"30",		-- 00e138: 3041             RET     
						   57657 => x"61",
						   -- Begin: __TI_decompress_none
						   57658 => x"0F",		-- 00e13a: 0F4C             MOV.W   R12,R15
						   57659 => x"6C",
						   57660 => x"0C",		-- 00e13c: 0C4D             MOV.W   R13,R12
						   57661 => x"6D",
						   57662 => x"3D",		-- 00e13e: 3D40             MOV.W   #0x0003,R13
						   57663 => x"60",
						   57664 => x"03",		-- 00e140: 0300            
						   57665 => x"00",
						   57666 => x"0D",		-- 00e142: 0D5F             ADD.W   R15,R13
						   57667 => x"7F",
						   57668 => x"1E",		-- 00e144: 1E4F             MOV.W   0x0001(R15),R14
						   57669 => x"6F",
						   57670 => x"01",		-- 00e146: 0100            
						   57671 => x"00",
						   57672 => x"30",		-- 00e148: 3040             BR      #memcpy
						   57673 => x"60",
						   57674 => x"5E",		-- 00e14a: 5EE1            
						   57675 => x"E1",
						   -- Begin: __mspabi_srll
						   57676 => x"3E",		-- 00e14c: 3EF0             AND.W   #0x001f,R14
						   57677 => x"10",
						   57678 => x"1F",		-- 00e14e: 1F00            
						   57679 => x"00",
						   57680 => x"05",		-- 00e150: 0524             JEQ     (L_LSR_RET)
						   57681 => x"44",
						   -- Begin: L_LSR_TOP
						   57682 => x"12",		-- 00e152: 12C3             CLRC    
						   57683 => x"E3",
						   57684 => x"0D",		-- 00e154: 0D10             RRC     R13
						   57685 => x"30",
						   57686 => x"0C",		-- 00e156: 0C10             RRC     R12
						   57687 => x"30",
						   57688 => x"1E",		-- 00e158: 1E83             DEC.W   R14
						   57689 => x"A3",
						   57690 => x"FB",		-- 00e15a: FB23             JNE     (L_LSR_TOP)
						   57691 => x"43",
						   -- Begin: L_LSR_RET
						   57692 => x"30",		-- 00e15c: 3041             RET     
						   57693 => x"61",
						   -- Begin: memcpy
						   57694 => x"0E",		-- 00e15e: 0E93             TST.W   R14
						   57695 => x"B3",
						   57696 => x"06",		-- 00e160: 0624             JEQ     ($C$L2)
						   57697 => x"44",
						   57698 => x"0F",		-- 00e162: 0F4C             MOV.W   R12,R15
						   57699 => x"6C",
						   57700 => x"1F",		-- 00e164: 1F53             INC.W   R15
						   57701 => x"73",
						   57702 => x"FF",		-- 00e166: FF4D             MOV.B   @R13+,0xffff(R15)
						   57703 => x"6D",
						   57704 => x"FF",		-- 00e168: FFFF            
						   57705 => x"FF",
						   57706 => x"1E",		-- 00e16a: 1E83             DEC.W   R14
						   57707 => x"A3",
						   57708 => x"FB",		-- 00e16c: FB23             JNE     ($C$L1)
						   57709 => x"43",
						   57710 => x"30",		-- 00e16e: 3041             RET     
						   57711 => x"61",
						   -- Begin: __mspabi_func_epilog_7
						   -- Begin: __mspabi_func_epilog
						   57712 => x"34",		-- 00e170: 3441             POP.W   R4
						   57713 => x"61",
						   -- Begin: __mspabi_func_epilog_6
						   57714 => x"35",		-- 00e172: 3541             POP.W   R5
						   57715 => x"61",
						   -- Begin: __mspabi_func_epilog_5
						   57716 => x"36",		-- 00e174: 3641             POP.W   R6
						   57717 => x"61",
						   -- Begin: __mspabi_func_epilog_4
						   57718 => x"37",		-- 00e176: 3741             POP.W   R7
						   57719 => x"61",
						   -- Begin: __mspabi_func_epilog_3
						   57720 => x"38",		-- 00e178: 3841             POP.W   R8
						   57721 => x"61",
						   -- Begin: __mspabi_func_epilog_2
						   57722 => x"39",		-- 00e17a: 3941             POP.W   R9
						   57723 => x"61",
						   -- Begin: __mspabi_func_epilog_1
						   57724 => x"3A",		-- 00e17c: 3A41             POP.W   R10
						   57725 => x"61",
						   57726 => x"30",		-- 00e17e: 3041             RET     
						   57727 => x"61",
						   -- Begin: strcpy
						   57728 => x"0F",		-- 00e180: 0F4C             MOV.W   R12,R15
						   57729 => x"6C",
						   57730 => x"7E",		-- 00e182: 7E4D             MOV.B   @R13+,R14
						   57731 => x"6D",
						   57732 => x"1F",		-- 00e184: 1F53             INC.W   R15
						   57733 => x"73",
						   57734 => x"CF",		-- 00e186: CF4E             MOV.B   R14,0xffff(R15)
						   57735 => x"6E",
						   57736 => x"FF",		-- 00e188: FFFF            
						   57737 => x"FF",
						   57738 => x"0E",		-- 00e18a: 0E93             TST.W   R14
						   57739 => x"B3",
						   57740 => x"FA",		-- 00e18c: FA23             JNE     ($C$L1)
						   57741 => x"43",
						   57742 => x"30",		-- 00e18e: 3041             RET     
						   57743 => x"61",
						   -- Begin: strlen
						   57744 => x"3F",		-- 00e190: 3F43             MOV.W   #-1,R15
						   57745 => x"63",
						   57746 => x"1F",		-- 00e192: 1F53             INC.W   R15
						   57747 => x"73",
						   57748 => x"7E",		-- 00e194: 7E4C             MOV.B   @R12+,R14
						   57749 => x"6C",
						   57750 => x"0E",		-- 00e196: 0E93             TST.W   R14
						   57751 => x"B3",
						   57752 => x"FC",		-- 00e198: FC23             JNE     ($C$L1)
						   57753 => x"43",
						   57754 => x"0C",		-- 00e19a: 0C4F             MOV.W   R15,R12
						   57755 => x"6F",
						   57756 => x"30",		-- 00e19c: 3041             RET     
						   57757 => x"61",
						   -- Begin: __mspabi_fltid
						   57758 => x"3C",		-- 00e19e: 3CB0             BIT.W   #0x8000,R12
						   57759 => x"D0",
						   57760 => x"00",		-- 00e1a0: 0080            
						   57761 => x"80",
						   57762 => x"0D",		-- 00e1a2: 0D7D             SUBC.W  R13,R13
						   57763 => x"9D",
						   57764 => x"3D",		-- 00e1a4: 3DE3             INV.W   R13
						   57765 => x"03",
						   57766 => x"30",		-- 00e1a6: 3040             BR      #__mspabi_fltlid
						   57767 => x"60",
						   57768 => x"A4",		-- 00e1a8: A4CE            
						   57769 => x"CE",
						   -- Begin: toupper
						   57770 => x"EC",		-- 00e1aa: ECB3             BIT.B   #2,0x992f(R12)
						   57771 => x"D3",
						   57772 => x"2F",		-- 00e1ac: 2F99            
						   57773 => x"99",
						   57774 => x"02",		-- 00e1ae: 0224             JEQ     ($C$L1)
						   57775 => x"44",
						   57776 => x"3C",		-- 00e1b0: 3C80             SUB.W   #0x0020,R12
						   57777 => x"A0",
						   57778 => x"20",		-- 00e1b2: 2000            
						   57779 => x"00",
						   57780 => x"30",		-- 00e1b4: 3041             RET     
						   57781 => x"61",
						   -- Begin: abs
						   57782 => x"0C",		-- 00e1b6: 0C93             TST.W   R12
						   57783 => x"B3",
						   57784 => x"02",		-- 00e1b8: 0234             JGE     ($C$L1)
						   57785 => x"54",
						   57786 => x"3C",		-- 00e1ba: 3CE3             INV.W   R12
						   57787 => x"03",
						   57788 => x"1C",		-- 00e1bc: 1C53             INC.W   R12
						   57789 => x"73",
						   57790 => x"30",		-- 00e1be: 3041             RET     
						   57791 => x"61",
						   -- Begin: malloc
						   57792 => x"0D",		-- 00e1c0: 0D4C             MOV.W   R12,R13
						   57793 => x"6C",
						   57794 => x"2C",		-- 00e1c2: 2C42             MOV.W   #4,R12
						   57795 => x"62",
						   57796 => x"30",		-- 00e1c4: 3040             BR      #aligned_alloc
						   57797 => x"60",
						   57798 => x"F2",		-- 00e1c6: F2C7            
						   57799 => x"C7",
						   -- Begin: _outc
						   57800 => x"4C",		-- 00e1c8: 4C4C             MOV.B   R12,R12
						   57801 => x"6C",
						   57802 => x"30",		-- 00e1ca: 3040             BR      #fputc
						   57803 => x"60",
						   57804 => x"8E",		-- 00e1cc: 8ED0            
						   57805 => x"D0",
						   -- Begin: abort
						   57806 => x"03",		-- 00e1ce: 0343             NOP     
						   57807 => x"63",
						   57808 => x"FF",		-- 00e1d0: FF3F             JMP     ($C$L1)
						   57809 => x"5F",
						   57810 => x"03",		-- 00e1d2: 0343             NOP     
						   57811 => x"63",
						   -- Begin: _outs
						   57812 => x"30",		-- 00e1d4: 3040             BR      #fputs
						   57813 => x"60",
						   57814 => x"E8",		-- 00e1d6: E8C8            
						   57815 => x"C8",
						   -- Begin: _system_pre_init
						   57816 => x"1C",		-- 00e1d8: 1C43             MOV.W   #1,R12
						   57817 => x"63",
						   57818 => x"30",		-- 00e1da: 3041             RET     
						   57819 => x"61",
						   -- Begin: _nop
						   57820 => x"30",		-- 00e1dc: 3041             RET     
						   57821 => x"61",
						   -- Begin: _system_post_cinit
						   57822 => x"30",		-- 00e1de: 3041             RET     
						   57823 => x"61",
						   -- ISR Trap
						   57824 => x"32",		-- 00e1e0: 32D0             BIS.W   #0x0010,SR
						   57825 => x"F0",
						   57826 => x"10",		-- 00e1e2: 1000            
						   57827 => x"00",
						   57828 => x"FD",		-- 00e1e4: FD3F             JMP     (__TI_ISR_TRAP)
						   57829 => x"5F",
						   57830 => x"03",		-- 00e1e6: 0343             NOP     
						   57831 => x"63",
						   -- IRQ Vectors (Interrupt Vectors)
						   65486 => x"e0",		-- 00ffce:e1e0 PORT4 __TI_int22 int22
						   65487 => x"e1",
						   65488 => x"e0",		-- 00ffd0:e1e0 PORT3 __TI_int23 int23
						   65489 => x"e1",
						   65490 => x"e0",		-- 00ffd2:e1e0 PORT2 __TI_int24 int24
						   65491 => x"e1",
						   65492 => x"e0",		-- 00ffd4:e1e0 PORT1 __TI_int25 int25
						   65493 => x"e1",
						   65494 => x"e0",		-- 00ffd6:e1e0 SAC1_SAC3 __TI_int26 int26
						   65495 => x"e1",
						   65496 => x"e0",		-- 00ffd8:e1e0 SAC0_SAC2 __TI_int27 int27
						   65497 => x"e1",
						   65498 => x"e0",		-- 00ffda:e1e0 ECOMP0_ECOMP1 __TI_int28 int28
						   65499 => x"e1",
						   65500 => x"e0",		-- 00ffdc:e1e0 ADC __TI_int29 int29
						   65501 => x"e1",
						   65502 => x"e0",		-- 00ffde:e1e0 EUSCI_B1 __TI_int30 int30
						   65503 => x"e1",
						   65504 => x"e0",		-- 00ffe0:e1e0 EUSCI_B0 __TI_int31 int31
						   65505 => x"e1",
						   65506 => x"e0",		-- 00ffe2:e1e0 EUSCI_A1 __TI_int32 int32
						   65507 => x"e1",
						   65508 => x"e0",		-- 00ffe4:e1e0 EUSCI_A0 __TI_int33 int33
						   65509 => x"e1",
						   65510 => x"e0",		-- 00ffe6:e1e0 WDT __TI_int34 int34
						   65511 => x"e1",
						   65512 => x"e0",		-- 00ffe8:e1e0 RTC __TI_int35 int35
						   65513 => x"e1",
						   65514 => x"e0",		-- 00ffea:e1e0 TIMER3_B1 __TI_int36 int36
						   65515 => x"e1",
						   65516 => x"e0",		-- 00ffec:e1e0 TIMER3_B0 __TI_int37 int37
						   65517 => x"e1",
						   65518 => x"e0",		-- 00ffee:e1e0 TIMER2_B1 __TI_int38 int38
						   65519 => x"e1",
						   65520 => x"e0",		-- 00fff0:e1e0 TIMER2_B0 __TI_int39 int39
						   65521 => x"e1",
						   65522 => x"e0",		-- 00fff2:e1e0 TIMER1_B1 __TI_int40 int40
						   65523 => x"e1",
						   65524 => x"e0",		-- 00fff4:e1e0 TIMER1_B0 __TI_int41 int41
						   65525 => x"e1",
						   65526 => x"e0",		-- 00fff6:e1e0 TIMER0_B1 __TI_int42 int42
						   65527 => x"e1",
						   65528 => x"e0",		-- 00fff8:e1e0 TIMER0_B0 __TI_int43 int43
						   65529 => x"e1",
						   65530 => x"e0",		-- 00fffa:e1e0 UNMI __TI_int44 int44
						   65531 => x"e1",
						   65532 => x"e0",		-- 00fffc:e1e0 SYSNMI __TI_int45 int45
						   65533 => x"e1",
						   65534 => x"44",		-- 00fffe:e044 .reset _reset_vector reset
						   65535 => x"e0",
						   others => x"00");

    signal EN : std_logic;
    
    begin
    -- Note 1:  The bus system uses a 16-bit Address (MAB)
    --          This address size can access locations from x0000 to xFFFF
    --          But our array is only defined from x8000 to xFFFF and
    --          if we try to access it with any other address, it will crash.
    --          So the first thing we need to do is create a local enable that
    --          will only assert when MAB is within x8000 to xFFFF.

     LOCAL_EN : process (MAB) 
     begin
         if ( (to_integer(unsigned(MAB)) >= 32768) and (to_integer(unsigned(MAB)) <= 65535)) then
           EN <= '1';
         else 
           EN <= '0';
         end if;
     end process;

    
    -- Note 2:  The bus system uses a 16-bit Address (MAB)
    --          The MDB_out is also provided as a 16-bit word
    --          However, the memory array is actually built as 8-bit bytes.
    --          So for a given 16-bit MAB, we give MDB_out = HB : LB
    --                                                 or  = ROM(MAB);1) : ROM(MAB)

    MEMORY_ROM : process (clk) 
    begin
        if (rising_edge(clk)) then
            if (EN='1' and write='0') then
                if(Byte = '0') then                      
                    MDB_in <= ROM(to_integer(unsigned(MAB)) + 1 ) & ROM(to_integer(unsigned(MAB)));
                else
                    MDB_in <= x"00" & ROM(to_integer(unsigned(MAB)));
                end if;
            end if;
        end if;
    end process;


end architecture;