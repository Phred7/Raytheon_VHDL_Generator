library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;


entity lowlife_memory is
    port ( clk	: in	std_logic;
         MAB		: in	std_logic_vector(15 downto 0);
         MDB_out  	: out	std_logic_vector(15 downto 0));
end entity;

architecture lowlife_memory_arch of lowlife_memory is

type rom_type is array (32768 to 65535) of std_logic_vector(7 downto 0);  -- this is MAB: x8000 to xFFFF
    
shared variable ROM : rom_type :=(32768 => x"00",		-- Begin: .cinit DATA Section
						   32769 => x"ff",
						   32770 => x"00",
						   32771 => x"38",
						   32772 => x"28",
						   32773 => x"37",
						   32774 => x"18",
						   32775 => x"00",
						   32776 => x"27",
						   32777 => x"34",
						   32778 => x"ff",
						   32779 => x"08",
						   32780 => x"39",
						   32781 => x"00",
						   32782 => x"00",
						   32783 => x"17",
						   32784 => x"00",
						   32785 => x"24",
						   32786 => x"0d",
						   32787 => x"ff",
						   32788 => x"78",
						   32789 => x"00",
						   32790 => x"29",
						   32791 => x"36",
						   32794 => x"00",
						   32795 => x"35",
						   32796 => x"fd",
						   32797 => x"07",
						   32798 => x"00",
						   32799 => x"40",
						   32800 => x"14",
						   32801 => x"13",
						   32802 => x"7d",
						   32803 => x"12",
						   32804 => x"68",
						   32805 => x"69",
						   32806 => x"ff",
						   32807 => x"00",
						   32808 => x"00",
						   32809 => x"19",
						   32810 => x"6a",
						   32811 => x"26",
						   32814 => x"3a",
						   32815 => x"be",
						   32816 => x"01",
						   32817 => x"50",
						   32818 => x"00",
						   32819 => x"25",
						   32820 => x"0e",
						   32821 => x"77",
						   32822 => x"76",
						   32823 => x"01",
						   32824 => x"d0",
						   32825 => x"6b",
						   32826 => x"ff",
						   32827 => x"00",
						   32828 => x"00",
						   32829 => x"04",
						   32830 => x"00",
						   32831 => x"03",
						   32832 => x"00",
						   32833 => x"6d",
						   32834 => x"6c",
						   32835 => x"df",
						   32836 => x"02",
						   32837 => x"01",
						   32838 => x"58",
						   32839 => x"00",
						   32840 => x"59",
						   32841 => x"01",
						   32842 => x"81",
						   32843 => x"33",
						   32844 => x"09",
						   32845 => x"ff",
						   32846 => x"0a",
						   32847 => x"5a",
						   32848 => x"00",
						   32849 => x"16",
						   32850 => x"0b",
						   32851 => x"00",
						   32852 => x"0c",
						   32853 => x"00",
						   32854 => x"e7",
						   32855 => x"00",
						   32856 => x"2a",
						   32857 => x"2b",
						   32858 => x"02",
						   32859 => x"91",
						   32860 => x"02",
						   32861 => x"d1",
						   32862 => x"15",
						   32863 => x"00",
						   32864 => x"7e",
						   32865 => x"af",
						   32866 => x"7f",
						   32867 => x"67",
						   32868 => x"00",
						   32869 => x"66",
						   32870 => x"00",
						   32871 => x"e4",
						   32872 => x"5b",
						   32873 => x"01",
						   32874 => x"62",
						   32875 => x"74",
						   32876 => x"ef",
						   32877 => x"75",
						   32880 => x"73",
						   32881 => x"06",
						   32882 => x"00",
						   32883 => x"5d",
						   32884 => x"5e",
						   32885 => x"5c",
						   32886 => x"ff",
						   32887 => x"00",
						   32888 => x"72",
						   32889 => x"5f",
						   32890 => x"71",
						   32891 => x"00",
						   32892 => x"48",
						   32893 => x"47",
						   32894 => x"00",
						   32895 => x"ff",
						   32896 => x"44",
						   32897 => x"49",
						   32900 => x"1d",
						   32901 => x"00",
						   32902 => x"46",
						   32903 => x"00",
						   32904 => x"ff",
						   32905 => x"45",
						   32908 => x"23",
						   32909 => x"22",
						   32910 => x"79",
						   32911 => x"00",
						   32912 => x"7a",
						   32913 => x"ff",
						   32914 => x"00",
						   32915 => x"4a",
						   32918 => x"1e",
						   32919 => x"06",
						   32920 => x"00",
						   32921 => x"7b",
						   32922 => x"f6",
						   32923 => x"08",
						   32924 => x"60",
						   32925 => x"7c",
						   32926 => x"11",
						   32927 => x"08",
						   32928 => x"b0",
						   32929 => x"43",
						   32930 => x"1a",
						   32931 => x"00",
						   32932 => x"1b",
						   32933 => x"57",
						   32934 => x"1c",
						   32935 => x"00",
						   32936 => x"3b",
						   32937 => x"05",
						   32938 => x"52",
						   32939 => x"0f",
						   32940 => x"05",
						   32941 => x"b5",
						   32942 => x"05",
						   32943 => x"0a",
						   32944 => x"40",
						   32945 => x"ff",
						   32946 => x"6e",
						   32947 => x"00",
						   32948 => x"6f",
						   32949 => x"10",
						   32950 => x"57",
						   32951 => x"54",
						   32952 => x"00",
						   32953 => x"2d",
						   32954 => x"af",
						   32955 => x"56",
						   32956 => x"55",
						   32957 => x"00",
						   32958 => x"32",
						   32959 => x"0b",
						   32960 => x"30",
						   32961 => x"2e",
						   32962 => x"0b",
						   32963 => x"70",
						   32964 => x"21",
						   32965 => x"ff",
						   32966 => x"00",
						   32967 => x"53",
						   32968 => x"00",
						   32969 => x"2c",
						   32970 => x"4b",
						   32971 => x"00",
						   32972 => x"00",
						   32973 => x"1f",
						   32974 => x"fe",
						   32975 => x"08",
						   32976 => x"34",
						   32977 => x"20",
						   32978 => x"64",
						   32979 => x"3d",
						   32980 => x"65",
						   32981 => x"42",
						   32982 => x"00",
						   32983 => x"3e",
						   32984 => x"bf",
						   32985 => x"00",
						   32986 => x"31",
						   32987 => x"63",
						   32988 => x"3c",
						   32989 => x"00",
						   32990 => x"2f",
						   32991 => x"0d",
						   32992 => x"70",
						   32993 => x"30",
						   32994 => x"ff",
						   32995 => x"4d",
						   32996 => x"52",
						   32997 => x"4e",
						   32998 => x"41",
						   32999 => x"4c",
						   33000 => x"3f",
						   33001 => x"00",
						   33002 => x"40",
						   33003 => x"ff",
						   33004 => x"62",
						   33005 => x"51",
						   33006 => x"4f",
						   33007 => x"50",
						   33008 => x"61",
						   33009 => x"60",
						   33010 => x"70",
						   33011 => x"00",
						   33012 => x"0f",
						   33013 => x"e8",
						   33014 => x"03",
						   33015 => x"3d",
						   33016 => x"00",
						   33017 => x"ff",
						   33018 => x"f0",
						   33019 => x"00",
						   33020 => x"c2",
						   33021 => x"81",
						   33022 => x"26",
						   33023 => x"83",
						   33024 => x"00",
						   33025 => x"80",
						   33026 => x"00",
						   33027 => x"20",
						   -- Begin: program memory TEXT Section
						   33028 => x"21",		-- 008104: 2183             DECD.W  SP
						   33029 => x"63",
						   33030 => x"B2",		-- 008106: B240             MOV.W   #0x5a80,&WDTCTL_L
						   33031 => x"20",
						   33032 => x"80",		-- 008108: 805A            
						   33033 => x"5A",
						   33034 => x"CC",		-- 00810a: CC01            
						   33035 => x"01",
						   33036 => x"92",		-- 00810c: 92C3             BIC.W   #1,&PM5CTL0_L
						   33037 => x"A3",
						   33038 => x"30",		-- 00810e: 3001            
						   33039 => x"01",
						   33040 => x"5F",		-- 008110: 5F42             MOV.B   &P1DIR,R15
						   33041 => x"22",
						   33042 => x"04",		-- 008112: 0402            
						   33043 => x"02",
						   33044 => x"C2",		-- 008114: C243             CLR.B   &P1DIR
						   33045 => x"23",
						   33046 => x"04",		-- 008116: 0402            
						   33047 => x"02",
						   33048 => x"F2",		-- 008118: F2F0             AND.B   #0x00fc,&P2DIR
						   33049 => x"D0",
						   33050 => x"FC",		-- 00811a: FC00            
						   33051 => x"00",
						   33052 => x"05",		-- 00811c: 0502            
						   33053 => x"02",
						   33054 => x"F2",		-- 00811e: F2D0             BIS.B   #0x0034,&P2DIR
						   33055 => x"B0",
						   33056 => x"34",		-- 008120: 3400            
						   33057 => x"00",
						   33058 => x"05",		-- 008122: 0502            
						   33059 => x"02",
						   33060 => x"B2",		-- 008124: B2D0             BIS.W   #0x0220,&TB0CTL_L
						   33061 => x"B0",
						   33062 => x"20",		-- 008126: 2002            
						   33063 => x"02",
						   33064 => x"80",		-- 008128: 8003            
						   33065 => x"03",
						   33066 => x"B2",		-- 00812a: B2D0             BIS.W   #0x0010,&TB0CCTL0_L
						   33067 => x"B0",
						   33068 => x"10",		-- 00812c: 1000            
						   33069 => x"00",
						   33070 => x"82",		-- 00812e: 8203            
						   33071 => x"03",
						   33072 => x"92",		-- 008130: 9242             MOV.W   &frequency,&TB0CCR0_L
						   33073 => x"22",
						   33074 => x"00",		-- 008132: 0021            
						   33075 => x"21",
						   33076 => x"92",		-- 008134: 9203            
						   33077 => x"03",
						   33078 => x"32",		-- 008136: 32D2             EINT    
						   33079 => x"B2",
						   33080 => x"3F",		-- 008138: 3F40             MOV.W   #0x0003,R15
						   33081 => x"20",
						   33082 => x"03",		-- 00813a: 0300            
						   33083 => x"00",
						   33084 => x"5F",		-- 00813c: 5FF2             AND.B   &P2IN,R15
						   33085 => x"D2",
						   33086 => x"01",		-- 00813e: 0102            
						   33087 => x"02",
						   33088 => x"C1",		-- 008140: C14F             MOV.B   R15,0x0000(SP)
						   33089 => x"2F",
						   33090 => x"00",		-- 008142: 0000            
						   33091 => x"00",
						   33092 => x"D1",		-- 008144: D193             CMP.B   #1,0x0000(SP)
						   33093 => x"73",
						   33094 => x"00",		-- 008146: 0000            
						   33095 => x"00",
						   33096 => x"04",		-- 008148: 0420             JNE     ($C$L2)
						   33097 => x"00",
						   33098 => x"B2",		-- 00814a: B240             MOV.W   #0x002f,&set_angle
						   33099 => x"20",
						   33100 => x"2F",		-- 00814c: 2F00            
						   33101 => x"00",
						   33102 => x"02",		-- 00814e: 0221            
						   33103 => x"21",
						   33104 => x"0A",		-- 008150: 0A3C             JMP     ($C$L4)
						   33105 => x"1C",
						   33106 => x"E1",		-- 008152: E193             CMP.B   #2,0x0000(SP)
						   33107 => x"73",
						   33108 => x"00",		-- 008154: 0000            
						   33109 => x"00",
						   33110 => x"04",		-- 008156: 0420             JNE     ($C$L3)
						   33111 => x"00",
						   33112 => x"B2",		-- 008158: B240             MOV.W   #0x004f,&set_angle
						   33113 => x"20",
						   33114 => x"4F",		-- 00815a: 4F00            
						   33115 => x"00",
						   33116 => x"02",		-- 00815c: 0221            
						   33117 => x"21",
						   33118 => x"03",		-- 00815e: 033C             JMP     ($C$L4)
						   33119 => x"1C",
						   33120 => x"B2",		-- 008160: B240             MOV.W   #0x003d,&set_angle
						   33121 => x"20",
						   33122 => x"3D",		-- 008162: 3D00            
						   33123 => x"00",
						   33124 => x"02",		-- 008164: 0221            
						   33125 => x"21",
						   33126 => x"5F",		-- 008166: 5F42             MOV.B   &P1IN,R15
						   33127 => x"22",
						   33128 => x"00",		-- 008168: 0002            
						   33129 => x"02",
						   33130 => x"D1",		-- 00816a: D14F             MOV.B   0x2000(R15),0x0000(SP)
						   33131 => x"2F",
						   33132 => x"00",		-- 00816c: 0020            
						   33133 => x"20",
						   33134 => x"00",		-- 00816e: 0000            
						   33135 => x"00",
						   33136 => x"6F",		-- 008170: 6F41             MOV.B   @SP,R15
						   33137 => x"21",
						   33138 => x"1F",		-- 008172: 1F92             CMP.W   &set_angle,R15
						   33139 => x"72",
						   33140 => x"02",		-- 008174: 0221            
						   33141 => x"21",
						   33142 => x"0B",		-- 008176: 0B2C             JHS     ($C$L5)
						   33143 => x"0C",
						   33144 => x"E2",		-- 008178: E2C2             BIC.B   #4,&P2OUT
						   33145 => x"A2",
						   33146 => x"03",		-- 00817a: 0302            
						   33147 => x"02",
						   33148 => x"F2",		-- 00817c: F2F0             AND.B   #0x00df,&P2OUT
						   33149 => x"D0",
						   33150 => x"DF",		-- 00817e: DF00            
						   33151 => x"00",
						   33152 => x"03",		-- 008180: 0302            
						   33153 => x"02",
						   33154 => x"5F",		-- 008182: 5F42             MOV.B   &set_angle,R15
						   33155 => x"22",
						   33156 => x"02",		-- 008184: 0221            
						   33157 => x"21",
						   33158 => x"6F",		-- 008186: 6F81             SUB.B   @SP,R15
						   33159 => x"61",
						   33160 => x"C1",		-- 008188: C14F             MOV.B   R15,0x0000(SP)
						   33161 => x"2F",
						   33162 => x"00",		-- 00818a: 0000            
						   33163 => x"00",
						   33164 => x"0F",		-- 00818c: 0F3C             JMP     ($C$L7)
						   33165 => x"1C",
						   33166 => x"6F",		-- 00818e: 6F41             MOV.B   @SP,R15
						   33167 => x"21",
						   33168 => x"82",		-- 008190: 829F             CMP.W   R15,&set_angle
						   33169 => x"7F",
						   33170 => x"02",		-- 008192: 0221            
						   33171 => x"21",
						   33172 => x"09",		-- 008194: 092C             JHS     ($C$L6)
						   33173 => x"0C",
						   33174 => x"E2",		-- 008196: E2C2             BIC.B   #4,&P2OUT
						   33175 => x"A2",
						   33176 => x"03",		-- 008198: 0302            
						   33177 => x"02",
						   33178 => x"F2",		-- 00819a: F2D0             BIS.B   #0x0020,&P2OUT
						   33179 => x"B0",
						   33180 => x"20",		-- 00819c: 2000            
						   33181 => x"00",
						   33182 => x"03",		-- 00819e: 0302            
						   33183 => x"02",
						   33184 => x"D1",		-- 0081a0: D182             SUB.B   &set_angle,0x0000(SP)
						   33185 => x"62",
						   33186 => x"02",		-- 0081a2: 0221            
						   33187 => x"21",
						   33188 => x"00",		-- 0081a4: 0000            
						   33189 => x"00",
						   33190 => x"02",		-- 0081a6: 023C             JMP     ($C$L7)
						   33191 => x"1C",
						   33192 => x"E2",		-- 0081a8: E2D2             BIS.B   #4,&P2OUT
						   33193 => x"B2",
						   33194 => x"03",		-- 0081aa: 0302            
						   33195 => x"02",
						   33196 => x"6F",		-- 0081ac: 6F41             MOV.B   @SP,R15
						   33197 => x"21",
						   33198 => x"0C",		-- 0081ae: 0C4F             MOV.W   R15,R12
						   33199 => x"2F",
						   33200 => x"B0",		-- 0081b0: B012             CALL    #__mspabi_slli_6
						   33201 => x"F2",
						   33202 => x"EA",		-- 0081b2: EA82            
						   33203 => x"82",
						   33204 => x"0C",		-- 0081b4: 0C8F             SUB.W   R15,R12
						   33205 => x"6F",
						   33206 => x"3F",		-- 0081b6: 3F40             MOV.W   #0x0fa0,R15
						   33207 => x"20",
						   33208 => x"A0",		-- 0081b8: A00F            
						   33209 => x"0F",
						   33210 => x"0F",		-- 0081ba: 0F8C             SUB.W   R12,R15
						   33211 => x"6C",
						   33212 => x"82",		-- 0081bc: 824F             MOV.W   R15,&frequency
						   33213 => x"2F",
						   33214 => x"00",		-- 0081be: 0021            
						   33215 => x"21",
						   33216 => x"BB",		-- 0081c0: BB3F             JMP     ($C$L1)
						   33217 => x"1F",
						   -- Begin: __TI_decompress_lzss
						   33218 => x"0A",		-- 0081c2: 0A12             PUSH    R10
						   33219 => x"F2",
						   33220 => x"09",		-- 0081c4: 0912             PUSH    R9
						   33221 => x"F2",
						   33222 => x"08",		-- 0081c6: 0812             PUSH    R8
						   33223 => x"F2",
						   33224 => x"0A",		-- 0081c8: 0A4C             MOV.W   R12,R10
						   33225 => x"2C",
						   33226 => x"78",		-- 0081ca: 784A             MOV.B   @R10+,R8
						   33227 => x"2A",
						   33228 => x"09",		-- 0081cc: 0943             CLR.W   R9
						   33229 => x"23",
						   33230 => x"11",		-- 0081ce: 113C             JMP     ($C$L6)
						   33231 => x"1C",
						   33232 => x"0E",		-- 0081d0: 0E4D             MOV.W   R13,R14
						   33233 => x"2D",
						   33234 => x"0E",		-- 0081d2: 0E8B             SUB.W   R11,R14
						   33235 => x"6B",
						   33236 => x"1E",		-- 0081d4: 1E83             DEC.W   R14
						   33237 => x"63",
						   33238 => x"1D",		-- 0081d6: 1D53             INC.W   R13
						   33239 => x"33",
						   33240 => x"FD",		-- 0081d8: FD4E             MOV.B   @R14+,0xffff(R13)
						   33241 => x"2E",
						   33242 => x"FF",		-- 0081da: FFFF            
						   33243 => x"FF",
						   33244 => x"1F",		-- 0081dc: 1F83             DEC.W   R15
						   33245 => x"63",
						   33246 => x"FB",		-- 0081de: FB23             JNE     ($C$L3)
						   33247 => x"03",
						   33248 => x"03",		-- 0081e0: 033C             JMP     ($C$L5)
						   33249 => x"1C",
						   33250 => x"1D",		-- 0081e2: 1D53             INC.W   R13
						   33251 => x"33",
						   33252 => x"FD",		-- 0081e4: FD4A             MOV.B   @R10+,0xffff(R13)
						   33253 => x"2A",
						   33254 => x"FF",		-- 0081e6: FFFF            
						   33255 => x"FF",
						   33256 => x"12",		-- 0081e8: 12C3             CLRC    
						   33257 => x"A3",
						   33258 => x"08",		-- 0081ea: 0810             RRC     R8
						   33259 => x"F0",
						   33260 => x"19",		-- 0081ec: 1953             INC.W   R9
						   33261 => x"33",
						   33262 => x"39",		-- 0081ee: 3992             CMP.W   #8,R9
						   33263 => x"72",
						   33264 => x"EC",		-- 0081f0: EC37             JGE     ($C$L1)
						   33265 => x"17",
						   33266 => x"18",		-- 0081f2: 18B3             BIT.W   #1,R8
						   33267 => x"93",
						   33268 => x"F6",		-- 0081f4: F623             JNE     ($C$L4)
						   33269 => x"03",
						   33270 => x"7B",		-- 0081f6: 7B4A             MOV.B   @R10+,R11
						   33271 => x"2A",
						   33272 => x"7F",		-- 0081f8: 7F4A             MOV.B   @R10+,R15
						   33273 => x"2A",
						   33274 => x"0C",		-- 0081fa: 0C4B             MOV.W   R11,R12
						   33275 => x"2B",
						   33276 => x"B0",		-- 0081fc: B012             CALL    #__mspabi_slli_4
						   33277 => x"F2",
						   33278 => x"EE",		-- 0081fe: EE82            
						   33279 => x"82",
						   33280 => x"0B",		-- 008200: 0B4C             MOV.W   R12,R11
						   33281 => x"2C",
						   33282 => x"0C",		-- 008202: 0C4F             MOV.W   R15,R12
						   33283 => x"2F",
						   33284 => x"B0",		-- 008204: B012             CALL    #__mspabi_srli_4
						   33285 => x"F2",
						   33286 => x"78",		-- 008206: 7882            
						   33287 => x"82",
						   33288 => x"3C",		-- 008208: 3CF0             AND.W   #0x000f,R12
						   33289 => x"D0",
						   33290 => x"0F",		-- 00820a: 0F00            
						   33291 => x"00",
						   33292 => x"0B",		-- 00820c: 0BDC             BIS.W   R12,R11
						   33293 => x"BC",
						   33294 => x"3F",		-- 00820e: 3FF0             AND.W   #0x000f,R15
						   33295 => x"D0",
						   33296 => x"0F",		-- 008210: 0F00            
						   33297 => x"00",
						   33298 => x"3F",		-- 008212: 3F50             ADD.W   #0x0003,R15
						   33299 => x"30",
						   33300 => x"03",		-- 008214: 0300            
						   33301 => x"00",
						   33302 => x"3F",		-- 008216: 3F90             CMP.W   #0x0012,R15
						   33303 => x"70",
						   33304 => x"12",		-- 008218: 1200            
						   33305 => x"00",
						   33306 => x"0C",		-- 00821a: 0C20             JNE     ($C$L8)
						   33307 => x"00",
						   33308 => x"7E",		-- 00821c: 7E4A             MOV.B   @R10+,R14
						   33309 => x"2A",
						   33310 => x"3E",		-- 00821e: 3EB0             BIT.W   #0x0080,R14
						   33311 => x"90",
						   33312 => x"80",		-- 008220: 8000            
						   33313 => x"00",
						   33314 => x"07",		-- 008222: 0724             JEQ     ($C$L7)
						   33315 => x"04",
						   33316 => x"7C",		-- 008224: 7C4A             MOV.B   @R10+,R12
						   33317 => x"2A",
						   33318 => x"4C",		-- 008226: 4C4C             MOV.B   R12,R12
						   33319 => x"2C",
						   33320 => x"B0",		-- 008228: B012             CALL    #__mspabi_slli_7
						   33321 => x"F2",
						   33322 => x"E8",		-- 00822a: E882            
						   33323 => x"82",
						   33324 => x"3E",		-- 00822c: 3EF0             AND.W   #0x007f,R14
						   33325 => x"D0",
						   33326 => x"7F",		-- 00822e: 7F00            
						   33327 => x"00",
						   33328 => x"0E",		-- 008230: 0EDC             BIS.W   R12,R14
						   33329 => x"BC",
						   33330 => x"0F",		-- 008232: 0F5E             ADD.W   R14,R15
						   33331 => x"3E",
						   33332 => x"3B",		-- 008234: 3B90             CMP.W   #0x0fff,R11
						   33333 => x"70",
						   33334 => x"FF",		-- 008236: FF0F            
						   33335 => x"0F",
						   33336 => x"CB",		-- 008238: CB23             JNE     ($C$L2)
						   33337 => x"03",
						   33338 => x"30",		-- 00823a: 3040             BR      #__mspabi_func_epilog_3
						   33339 => x"20",
						   33340 => x"52",		-- 00823c: 5283            
						   33341 => x"83",
						   -- Begin: __mspabi_srli
						   33342 => x"3D",		-- 00823e: 3DF0             AND.W   #0x000f,R13
						   33343 => x"D0",
						   33344 => x"0F",		-- 008240: 0F00            
						   33345 => x"00",
						   33346 => x"3D",		-- 008242: 3DE0             XOR.W   #0x000f,R13
						   33347 => x"C0",
						   33348 => x"0F",		-- 008244: 0F00            
						   33349 => x"00",
						   33350 => x"0D",		-- 008246: 0D5D             RLA.W   R13
						   33351 => x"3D",
						   33352 => x"0D",		-- 008248: 0D5D             RLA.W   R13
						   33353 => x"3D",
						   33354 => x"00",		-- 00824a: 005D             ADD.W   R13,PC
						   33355 => x"3D",
						   -- Begin: __mspabi_srli_15
						   33356 => x"12",		-- 00824c: 12C3             CLRC    
						   33357 => x"A3",
						   33358 => x"0C",		-- 00824e: 0C10             RRC     R12
						   33359 => x"F0",
						   -- Begin: __mspabi_srli_14
						   33360 => x"12",		-- 008250: 12C3             CLRC    
						   33361 => x"A3",
						   33362 => x"0C",		-- 008252: 0C10             RRC     R12
						   33363 => x"F0",
						   -- Begin: __mspabi_srli_13
						   33364 => x"12",		-- 008254: 12C3             CLRC    
						   33365 => x"A3",
						   33366 => x"0C",		-- 008256: 0C10             RRC     R12
						   33367 => x"F0",
						   -- Begin: __mspabi_srli_12
						   33368 => x"12",		-- 008258: 12C3             CLRC    
						   33369 => x"A3",
						   33370 => x"0C",		-- 00825a: 0C10             RRC     R12
						   33371 => x"F0",
						   -- Begin: __mspabi_srli_11
						   33372 => x"12",		-- 00825c: 12C3             CLRC    
						   33373 => x"A3",
						   33374 => x"0C",		-- 00825e: 0C10             RRC     R12
						   33375 => x"F0",
						   -- Begin: __mspabi_srli_10
						   33376 => x"12",		-- 008260: 12C3             CLRC    
						   33377 => x"A3",
						   33378 => x"0C",		-- 008262: 0C10             RRC     R12
						   33379 => x"F0",
						   -- Begin: __mspabi_srli_9
						   33380 => x"12",		-- 008264: 12C3             CLRC    
						   33381 => x"A3",
						   33382 => x"0C",		-- 008266: 0C10             RRC     R12
						   33383 => x"F0",
						   -- Begin: __mspabi_srli_8
						   33384 => x"12",		-- 008268: 12C3             CLRC    
						   33385 => x"A3",
						   33386 => x"0C",		-- 00826a: 0C10             RRC     R12
						   33387 => x"F0",
						   -- Begin: __mspabi_srli_7
						   33388 => x"12",		-- 00826c: 12C3             CLRC    
						   33389 => x"A3",
						   33390 => x"0C",		-- 00826e: 0C10             RRC     R12
						   33391 => x"F0",
						   -- Begin: __mspabi_srli_6
						   33392 => x"12",		-- 008270: 12C3             CLRC    
						   33393 => x"A3",
						   33394 => x"0C",		-- 008272: 0C10             RRC     R12
						   33395 => x"F0",
						   -- Begin: __mspabi_srli_5
						   33396 => x"12",		-- 008274: 12C3             CLRC    
						   33397 => x"A3",
						   33398 => x"0C",		-- 008276: 0C10             RRC     R12
						   33399 => x"F0",
						   -- Begin: __mspabi_srli_4
						   33400 => x"12",		-- 008278: 12C3             CLRC    
						   33401 => x"A3",
						   33402 => x"0C",		-- 00827a: 0C10             RRC     R12
						   33403 => x"F0",
						   -- Begin: __mspabi_srli_3
						   33404 => x"12",		-- 00827c: 12C3             CLRC    
						   33405 => x"A3",
						   33406 => x"0C",		-- 00827e: 0C10             RRC     R12
						   33407 => x"F0",
						   -- Begin: __mspabi_srli_2
						   33408 => x"12",		-- 008280: 12C3             CLRC    
						   33409 => x"A3",
						   33410 => x"0C",		-- 008282: 0C10             RRC     R12
						   33411 => x"F0",
						   -- Begin: __mspabi_srli_1
						   33412 => x"12",		-- 008284: 12C3             CLRC    
						   33413 => x"A3",
						   33414 => x"0C",		-- 008286: 0C10             RRC     R12
						   33415 => x"F0",
						   33416 => x"30",		-- 008288: 3041             RET     
						   33417 => x"21",
						   -- Begin: __TI_auto_init_nobinit_nopinit
						   33418 => x"0A",		-- 00828a: 0A12             PUSH    R10
						   33419 => x"F2",
						   33420 => x"09",		-- 00828c: 0912             PUSH    R9
						   33421 => x"F2",
						   33422 => x"3F",		-- 00828e: 3F40             MOV.W   #0x80fc,R15
						   33423 => x"20",
						   33424 => x"FC",		-- 008290: FC80            
						   33425 => x"80",
						   33426 => x"3F",		-- 008292: 3F90             CMP.W   #0x8100,R15
						   33427 => x"70",
						   33428 => x"00",		-- 008294: 0081            
						   33429 => x"81",
						   33430 => x"16",		-- 008296: 1624             JEQ     ($C$L22)
						   33431 => x"04",
						   33432 => x"3F",		-- 008298: 3F40             MOV.W   #0x8100,R15
						   33433 => x"20",
						   33434 => x"00",		-- 00829a: 0081            
						   33435 => x"81",
						   33436 => x"3F",		-- 00829c: 3F90             CMP.W   #0x8104,R15
						   33437 => x"70",
						   33438 => x"04",		-- 00829e: 0481            
						   33439 => x"81",
						   33440 => x"11",		-- 0082a0: 1124             JEQ     ($C$L22)
						   33441 => x"04",
						   33442 => x"3A",		-- 0082a2: 3A40             MOV.W   #0x8104,R10
						   33443 => x"20",
						   33444 => x"04",		-- 0082a4: 0481            
						   33445 => x"81",
						   33446 => x"3A",		-- 0082a6: 3A80             SUB.W   #0x8100,R10
						   33447 => x"60",
						   33448 => x"00",		-- 0082a8: 0081            
						   33449 => x"81",
						   33450 => x"0A",		-- 0082aa: 0A11             RRA     R10
						   33451 => x"F1",
						   33452 => x"0A",		-- 0082ac: 0A11             RRA     R10
						   33453 => x"F1",
						   33454 => x"39",		-- 0082ae: 3940             MOV.W   #0x8100,R9
						   33455 => x"20",
						   33456 => x"00",		-- 0082b0: 0081            
						   33457 => x"81",
						   33458 => x"3C",		-- 0082b2: 3C49             MOV.W   @R9+,R12
						   33459 => x"29",
						   33460 => x"7F",		-- 0082b4: 7F4C             MOV.B   @R12+,R15
						   33461 => x"2C",
						   33462 => x"0F",		-- 0082b6: 0F5F             RLA.W   R15
						   33463 => x"3F",
						   33464 => x"1F",		-- 0082b8: 1F4F             MOV.W   0x80fc(R15),R15
						   33465 => x"2F",
						   33466 => x"FC",		-- 0082ba: FC80            
						   33467 => x"80",
						   33468 => x"3D",		-- 0082bc: 3D49             MOV.W   @R9+,R13
						   33469 => x"29",
						   33470 => x"8F",		-- 0082be: 8F12             CALL    R15
						   33471 => x"F2",
						   33472 => x"1A",		-- 0082c0: 1A83             DEC.W   R10
						   33473 => x"63",
						   33474 => x"F7",		-- 0082c2: F723             JNE     ($C$L21)
						   33475 => x"03",
						   33476 => x"B0",		-- 0082c4: B012             CALL    #_system_post_cinit
						   33477 => x"F2",
						   33478 => x"64",		-- 0082c6: 6483            
						   33479 => x"83",
						   33480 => x"30",		-- 0082c8: 3040             BR      #__mspabi_func_epilog_2
						   33481 => x"20",
						   33482 => x"54",		-- 0082ca: 5483            
						   33483 => x"83",
						   -- Begin: __mspabi_slli
						   33484 => x"3D",		-- 0082cc: 3DF0             AND.W   #0x000f,R13
						   33485 => x"D0",
						   33486 => x"0F",		-- 0082ce: 0F00            
						   33487 => x"00",
						   33488 => x"3D",		-- 0082d0: 3DE0             XOR.W   #0x000f,R13
						   33489 => x"C0",
						   33490 => x"0F",		-- 0082d2: 0F00            
						   33491 => x"00",
						   33492 => x"0D",		-- 0082d4: 0D5D             RLA.W   R13
						   33493 => x"3D",
						   33494 => x"00",		-- 0082d6: 005D             ADD.W   R13,PC
						   33495 => x"3D",
						   -- Begin: __mspabi_slli_15
						   33496 => x"0C",		-- 0082d8: 0C5C             RLA.W   R12
						   33497 => x"3C",
						   -- Begin: __mspabi_slli_14
						   33498 => x"0C",		-- 0082da: 0C5C             RLA.W   R12
						   33499 => x"3C",
						   -- Begin: __mspabi_slli_13
						   33500 => x"0C",		-- 0082dc: 0C5C             RLA.W   R12
						   33501 => x"3C",
						   -- Begin: __mspabi_slli_12
						   33502 => x"0C",		-- 0082de: 0C5C             RLA.W   R12
						   33503 => x"3C",
						   -- Begin: __mspabi_slli_11
						   33504 => x"0C",		-- 0082e0: 0C5C             RLA.W   R12
						   33505 => x"3C",
						   -- Begin: __mspabi_slli_10
						   33506 => x"0C",		-- 0082e2: 0C5C             RLA.W   R12
						   33507 => x"3C",
						   -- Begin: __mspabi_slli_9
						   33508 => x"0C",		-- 0082e4: 0C5C             RLA.W   R12
						   33509 => x"3C",
						   -- Begin: __mspabi_slli_8
						   33510 => x"0C",		-- 0082e6: 0C5C             RLA.W   R12
						   33511 => x"3C",
						   -- Begin: __mspabi_slli_7
						   33512 => x"0C",		-- 0082e8: 0C5C             RLA.W   R12
						   33513 => x"3C",
						   -- Begin: __mspabi_slli_6
						   33514 => x"0C",		-- 0082ea: 0C5C             RLA.W   R12
						   33515 => x"3C",
						   -- Begin: __mspabi_slli_5
						   33516 => x"0C",		-- 0082ec: 0C5C             RLA.W   R12
						   33517 => x"3C",
						   -- Begin: __mspabi_slli_4
						   33518 => x"0C",		-- 0082ee: 0C5C             RLA.W   R12
						   33519 => x"3C",
						   -- Begin: __mspabi_slli_3
						   33520 => x"0C",		-- 0082f0: 0C5C             RLA.W   R12
						   33521 => x"3C",
						   -- Begin: __mspabi_slli_2
						   33522 => x"0C",		-- 0082f2: 0C5C             RLA.W   R12
						   33523 => x"3C",
						   -- Begin: __mspabi_slli_1
						   33524 => x"0C",		-- 0082f4: 0C5C             RLA.W   R12
						   33525 => x"3C",
						   33526 => x"30",		-- 0082f6: 3041             RET     
						   33527 => x"21",
						   -- Begin: _c_int00_noargs
						   33528 => x"31",		-- 0082f8: 3140             MOV.W   #0x3000,SP
						   33529 => x"20",
						   33530 => x"00",		-- 0082fa: 0030            
						   33531 => x"30",
						   33532 => x"B0",		-- 0082fc: B012             CALL    #_system_pre_init
						   33533 => x"F2",
						   33534 => x"60",		-- 0082fe: 6083            
						   33535 => x"83",
						   33536 => x"0C",		-- 008300: 0C93             TST.W   R12
						   33537 => x"73",
						   33538 => x"02",		-- 008302: 0224             JEQ     ($C$L2)
						   33539 => x"04",
						   33540 => x"B0",		-- 008304: B012             CALL    #__TI_auto_init_nobinit_nopinit
						   33541 => x"F2",
						   33542 => x"8A",		-- 008306: 8A82            
						   33543 => x"82",
						   33544 => x"0C",		-- 008308: 0C43             CLR.W   R12
						   33545 => x"23",
						   33546 => x"B0",		-- 00830a: B012             CALL    #main
						   33547 => x"F2",
						   33548 => x"04",		-- 00830c: 0481            
						   33549 => x"81",
						   33550 => x"1C",		-- 00830e: 1C43             MOV.W   #1,R12
						   33551 => x"23",
						   33552 => x"B0",		-- 008310: B012             CALL    #abort
						   33553 => x"F2",
						   33554 => x"5A",		-- 008312: 5A83            
						   33555 => x"83",
						   -- Begin: Timer_ISR
						   33556 => x"92",		-- 008314: 9252             ADD.W   &frequency,&TB0CCR0_L
						   33557 => x"32",
						   33558 => x"00",		-- 008316: 0021            
						   33559 => x"21",
						   33560 => x"92",		-- 008318: 9203            
						   33561 => x"03",
						   33562 => x"F2",		-- 00831a: F2E0             XOR.B   #0x0010,&P2OUT
						   33563 => x"C0",
						   33564 => x"10",		-- 00831c: 1000            
						   33565 => x"00",
						   33566 => x"03",		-- 00831e: 0302            
						   33567 => x"02",
						   33568 => x"92",		-- 008320: 92C3             BIC.W   #1,&TB0CCTL0_L
						   33569 => x"A3",
						   33570 => x"82",		-- 008322: 8203            
						   33571 => x"03",
						   33572 => x"00",		-- 008324: 0013             RETI    
						   33573 => x"F3",
						   -- Begin: __TI_decompress_none
						   33574 => x"0F",		-- 008326: 0F4C             MOV.W   R12,R15
						   33575 => x"2C",
						   33576 => x"0C",		-- 008328: 0C4D             MOV.W   R13,R12
						   33577 => x"2D",
						   33578 => x"3D",		-- 00832a: 3D40             MOV.W   #0x0003,R13
						   33579 => x"20",
						   33580 => x"03",		-- 00832c: 0300            
						   33581 => x"00",
						   33582 => x"0D",		-- 00832e: 0D5F             ADD.W   R15,R13
						   33583 => x"3F",
						   33584 => x"1E",		-- 008330: 1E4F             MOV.W   0x0001(R15),R14
						   33585 => x"2F",
						   33586 => x"01",		-- 008332: 0100            
						   33587 => x"00",
						   33588 => x"30",		-- 008334: 3040             BR      #memcpy
						   33589 => x"20",
						   33590 => x"38",		-- 008336: 3883            
						   33591 => x"83",
						   -- Begin: memcpy
						   33592 => x"0E",		-- 008338: 0E93             TST.W   R14
						   33593 => x"73",
						   33594 => x"06",		-- 00833a: 0624             JEQ     ($C$L2)
						   33595 => x"04",
						   33596 => x"0F",		-- 00833c: 0F4C             MOV.W   R12,R15
						   33597 => x"2C",
						   33598 => x"1F",		-- 00833e: 1F53             INC.W   R15
						   33599 => x"33",
						   33600 => x"FF",		-- 008340: FF4D             MOV.B   @R13+,0xffff(R15)
						   33601 => x"2D",
						   33602 => x"FF",		-- 008342: FFFF            
						   33603 => x"FF",
						   33604 => x"1E",		-- 008344: 1E83             DEC.W   R14
						   33605 => x"63",
						   33606 => x"FB",		-- 008346: FB23             JNE     ($C$L1)
						   33607 => x"03",
						   33608 => x"30",		-- 008348: 3041             RET     
						   33609 => x"21",
						   -- Begin: __mspabi_func_epilog_7
						   -- Begin: __mspabi_func_epilog
						   33610 => x"34",		-- 00834a: 3441             POP.W   R4
						   33611 => x"21",
						   -- Begin: __mspabi_func_epilog_6
						   33612 => x"35",		-- 00834c: 3541             POP.W   R5
						   33613 => x"21",
						   -- Begin: __mspabi_func_epilog_5
						   33614 => x"36",		-- 00834e: 3641             POP.W   R6
						   33615 => x"21",
						   -- Begin: __mspabi_func_epilog_4
						   33616 => x"37",		-- 008350: 3741             POP.W   R7
						   33617 => x"21",
						   -- Begin: __mspabi_func_epilog_3
						   33618 => x"38",		-- 008352: 3841             POP.W   R8
						   33619 => x"21",
						   -- Begin: __mspabi_func_epilog_2
						   33620 => x"39",		-- 008354: 3941             POP.W   R9
						   33621 => x"21",
						   -- Begin: __mspabi_func_epilog_1
						   33622 => x"3A",		-- 008356: 3A41             POP.W   R10
						   33623 => x"21",
						   33624 => x"30",		-- 008358: 3041             RET     
						   33625 => x"21",
						   -- Begin: abort
						   33626 => x"03",		-- 00835a: 0343             NOP     
						   33627 => x"23",
						   33628 => x"FF",		-- 00835c: FF3F             JMP     ($C$L1)
						   33629 => x"1F",
						   33630 => x"03",		-- 00835e: 0343             NOP     
						   33631 => x"23",
						   -- Begin: _system_pre_init
						   33632 => x"1C",		-- 008360: 1C43             MOV.W   #1,R12
						   33633 => x"23",
						   33634 => x"30",		-- 008362: 3041             RET     
						   33635 => x"21",
						   -- Begin: _system_post_cinit
						   33636 => x"30",		-- 008364: 3041             RET     
						   33637 => x"21",
						   -- ISR Trap
						   33638 => x"32",		-- 008366: 32D0             BIS.W   #0x0010,SR
						   33639 => x"B0",
						   33640 => x"10",		-- 008368: 1000            
						   33641 => x"00",
						   33642 => x"FD",		-- 00836a: FD3F             JMP     (__TI_ISR_TRAP)
						   33643 => x"1F",
						   33644 => x"03",		-- 00836c: 0343             NOP     
						   33645 => x"23",
						   -- IRQ Vectors (Interrupt Vectors)
						   65486 => x"66",		-- 00ffce:8366 PORT4 __TI_int22 int22
						   65487 => x"83",
						   65488 => x"66",		-- 00ffd0:8366 PORT3 __TI_int23 int23
						   65489 => x"83",
						   65490 => x"66",		-- 00ffd2:8366 PORT2 __TI_int24 int24
						   65491 => x"83",
						   65492 => x"66",		-- 00ffd4:8366 PORT1 __TI_int25 int25
						   65493 => x"83",
						   65494 => x"66",		-- 00ffd6:8366 SAC1_SAC3 __TI_int26 int26
						   65495 => x"83",
						   65496 => x"66",		-- 00ffd8:8366 SAC0_SAC2 __TI_int27 int27
						   65497 => x"83",
						   65498 => x"66",		-- 00ffda:8366 ECOMP0_ECOMP1 __TI_int28 int28
						   65499 => x"83",
						   65500 => x"66",		-- 00ffdc:8366 ADC __TI_int29 int29
						   65501 => x"83",
						   65502 => x"66",		-- 00ffde:8366 EUSCI_B1 __TI_int30 int30
						   65503 => x"83",
						   65504 => x"66",		-- 00ffe0:8366 EUSCI_B0 __TI_int31 int31
						   65505 => x"83",
						   65506 => x"66",		-- 00ffe2:8366 EUSCI_A1 __TI_int32 int32
						   65507 => x"83",
						   65508 => x"66",		-- 00ffe4:8366 EUSCI_A0 __TI_int33 int33
						   65509 => x"83",
						   65510 => x"66",		-- 00ffe6:8366 WDT __TI_int34 int34
						   65511 => x"83",
						   65512 => x"66",		-- 00ffe8:8366 RTC __TI_int35 int35
						   65513 => x"83",
						   65514 => x"66",		-- 00ffea:8366 TIMER3_B1 __TI_int36 int36
						   65515 => x"83",
						   65516 => x"66",		-- 00ffec:8366 TIMER3_B0 __TI_int37 int37
						   65517 => x"83",
						   65518 => x"66",		-- 00ffee:8366 TIMER2_B1 __TI_int38 int38
						   65519 => x"83",
						   65520 => x"66",		-- 00fff0:8366 TIMER2_B0 __TI_int39 int39
						   65521 => x"83",
						   65522 => x"66",		-- 00fff2:8366 TIMER1_B1 __TI_int40 int40
						   65523 => x"83",
						   65524 => x"66",		-- 00fff4:8366 TIMER1_B0 __TI_int41 int41
						   65525 => x"83",
						   65526 => x"66",		-- 00fff6:8366 TIMER0_B1 __TI_int42 int42
						   65527 => x"83",
						   65528 => x"14",		-- 00fff8:8314 TIMER0_B0 __TI_int43 int43
						   65529 => x"83",
						   65530 => x"66",		-- 00fffa:8366 UNMI __TI_int44 int44
						   65531 => x"83",
						   65532 => x"66",		-- 00fffc:8366 SYSNMI __TI_int45 int45
						   65533 => x"83",
						   65534 => x"f8",		-- 00fffe:82f8 .reset _reset_vector reset
						   65535 => x"82",
						   others => x"00");

    
    signal high_addr, low_addr : integer;
    signal read_value : std_logic_vector(15 downto 0);
    signal EN : std_logic;
        
    
    begin
    -- Note 1:  The bus system uses a 16-bit Address (MAB)
    --          This address size can access locations from x0000 to xFFFF
    --          But our array is only defined from x8000 to xFFFF and
    --          if we try to access it with any other address, it will crash.
    --          So the first thing we need to do is create a local enable that
    --          will only assert when MAB is within x8000 to xFFFF.
     LOCAL_EN : process (MAB) 
     begin
         if ( (to_integer(unsigned(MAB)) >= 32768) and (to_integer(unsigned(MAB)) <= 65535)) then
           EN <= '1';
         else 
           EN <= '0';
         end if;
     end process;
    -- Note 2:  The bus system uses a 16-bit Address (MAB)
    --          The MDB_out is also provided as a 16-bit word
    --          However, the memory array is actually built as 8-bit bytes.
    --          So for a given 16-bit MAB, we give MDB_out = HB : LB
    --                                                 or  = RW(MAB+1) : RW(MAB)
    ADDR_HANDLE : process( MAB )
    begin
        if ( (to_integer(unsigned(MAB)) >= 32768) and (to_integer(unsigned(MAB)) <= 65535)) then
            high_addr<= to_integer(unsigned(MAB))+1;
            low_addr<= to_integer(unsigned(MAB));
        else
            high_addr<= 32769;
            low_addr <= 32768;   
        end if;
    end process ; -- ADDR_HANDLE
    LOW_BYTE : process(clk) 
    begin
        if (rising_edge(clk)) then
            read_value(7 downto 0) <= ROM(low_addr);
        end if;
    end process ; -- LOW_BYTE
    WRITE_HIGH_BYTE : process( clk )
    begin
        if (rising_edge(clk)) then
            read_value(15 downto 8)<=ROM(high_addr);
        end if ;
    end process ; -- WRITE_HIGH_BYTE
    MDB_out <= read_value;
    --------------------------------------------------------------------------------------------

end architecture;