library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;


entity highroller_memory is
    port ( clk	: in	std_logic;
         MAB		: in	std_logic_vector(15 downto 0);
         MDB_in  	: out	std_logic_vector(15 downto 0);
         MDB_out  	: in	std_logic_vector(15 downto 0);
         write	    : in	std_logic;
         Byte       : in    std_logic);
end entity;

architecture highroller_memory_arch of highroller_memory is

type rom_type is array (32768 to 65535) of std_logic_vector(7 downto 0);  -- this is MAB: x8000 to xFFFF
    
constant ROM : rom_type :=(32768 => x"00",		-- Begin: .cinit DATA Section
						   32769 => x"ff",
						   32770 => x"00",
						   32771 => x"38",
						   32772 => x"28",
						   32773 => x"37",
						   32774 => x"18",
						   32775 => x"00",
						   32776 => x"27",
						   32777 => x"34",
						   32778 => x"ff",
						   32779 => x"08",
						   32780 => x"39",
						   32781 => x"00",
						   32782 => x"00",
						   32783 => x"17",
						   32784 => x"00",
						   32785 => x"24",
						   32786 => x"0d",
						   32787 => x"ff",
						   32788 => x"78",
						   32789 => x"00",
						   32790 => x"29",
						   32791 => x"36",
						   32794 => x"00",
						   32795 => x"35",
						   32796 => x"fd",
						   32797 => x"07",
						   32798 => x"00",
						   32799 => x"40",
						   32800 => x"14",
						   32801 => x"13",
						   32802 => x"7d",
						   32803 => x"12",
						   32804 => x"68",
						   32805 => x"69",
						   32806 => x"ff",
						   32807 => x"00",
						   32808 => x"00",
						   32809 => x"19",
						   32810 => x"6a",
						   32811 => x"26",
						   32814 => x"3a",
						   32815 => x"be",
						   32816 => x"01",
						   32817 => x"50",
						   32818 => x"00",
						   32819 => x"25",
						   32820 => x"0e",
						   32821 => x"77",
						   32822 => x"76",
						   32823 => x"01",
						   32824 => x"d0",
						   32825 => x"6b",
						   32826 => x"ff",
						   32827 => x"00",
						   32828 => x"00",
						   32829 => x"04",
						   32830 => x"00",
						   32831 => x"03",
						   32832 => x"00",
						   32833 => x"6d",
						   32834 => x"6c",
						   32835 => x"df",
						   32836 => x"02",
						   32837 => x"01",
						   32838 => x"58",
						   32839 => x"00",
						   32840 => x"59",
						   32841 => x"01",
						   32842 => x"81",
						   32843 => x"33",
						   32844 => x"09",
						   32845 => x"ff",
						   32846 => x"0a",
						   32847 => x"5a",
						   32848 => x"00",
						   32849 => x"16",
						   32850 => x"0b",
						   32851 => x"00",
						   32852 => x"0c",
						   32853 => x"00",
						   32854 => x"e7",
						   32855 => x"00",
						   32856 => x"2a",
						   32857 => x"2b",
						   32858 => x"02",
						   32859 => x"91",
						   32860 => x"02",
						   32861 => x"d1",
						   32862 => x"15",
						   32863 => x"00",
						   32864 => x"7e",
						   32865 => x"af",
						   32866 => x"7f",
						   32867 => x"67",
						   32868 => x"00",
						   32869 => x"66",
						   32870 => x"00",
						   32871 => x"e4",
						   32872 => x"5b",
						   32873 => x"01",
						   32874 => x"62",
						   32875 => x"74",
						   32876 => x"ef",
						   32877 => x"75",
						   32880 => x"73",
						   32881 => x"06",
						   32882 => x"00",
						   32883 => x"5d",
						   32884 => x"5e",
						   32885 => x"5c",
						   32886 => x"ff",
						   32887 => x"00",
						   32888 => x"72",
						   32889 => x"5f",
						   32890 => x"71",
						   32891 => x"00",
						   32892 => x"48",
						   32893 => x"47",
						   32894 => x"00",
						   32895 => x"ff",
						   32896 => x"44",
						   32897 => x"49",
						   32900 => x"1d",
						   32901 => x"00",
						   32902 => x"46",
						   32903 => x"00",
						   32904 => x"ff",
						   32905 => x"45",
						   32908 => x"23",
						   32909 => x"22",
						   32910 => x"79",
						   32911 => x"00",
						   32912 => x"7a",
						   32913 => x"ff",
						   32914 => x"00",
						   32915 => x"4a",
						   32918 => x"1e",
						   32919 => x"06",
						   32920 => x"00",
						   32921 => x"7b",
						   32922 => x"f6",
						   32923 => x"08",
						   32924 => x"60",
						   32925 => x"7c",
						   32926 => x"11",
						   32927 => x"08",
						   32928 => x"b0",
						   32929 => x"43",
						   32930 => x"1a",
						   32931 => x"00",
						   32932 => x"1b",
						   32933 => x"57",
						   32934 => x"1c",
						   32935 => x"00",
						   32936 => x"3b",
						   32937 => x"05",
						   32938 => x"52",
						   32939 => x"0f",
						   32940 => x"05",
						   32941 => x"b5",
						   32942 => x"05",
						   32943 => x"0a",
						   32944 => x"40",
						   32945 => x"ff",
						   32946 => x"6e",
						   32947 => x"00",
						   32948 => x"6f",
						   32949 => x"10",
						   32950 => x"57",
						   32951 => x"54",
						   32952 => x"00",
						   32953 => x"2d",
						   32954 => x"af",
						   32955 => x"56",
						   32956 => x"55",
						   32957 => x"00",
						   32958 => x"32",
						   32959 => x"0b",
						   32960 => x"30",
						   32961 => x"2e",
						   32962 => x"0b",
						   32963 => x"70",
						   32964 => x"21",
						   32965 => x"ff",
						   32966 => x"00",
						   32967 => x"53",
						   32968 => x"00",
						   32969 => x"2c",
						   32970 => x"4b",
						   32971 => x"00",
						   32972 => x"00",
						   32973 => x"1f",
						   32974 => x"fe",
						   32975 => x"08",
						   32976 => x"34",
						   32977 => x"20",
						   32978 => x"64",
						   32979 => x"3d",
						   32980 => x"65",
						   32981 => x"42",
						   32982 => x"00",
						   32983 => x"3e",
						   32984 => x"bf",
						   32985 => x"00",
						   32986 => x"31",
						   32987 => x"63",
						   32988 => x"3c",
						   32989 => x"00",
						   32990 => x"2f",
						   32991 => x"0d",
						   32992 => x"70",
						   32993 => x"30",
						   32994 => x"ff",
						   32995 => x"4d",
						   32996 => x"52",
						   32997 => x"4e",
						   32998 => x"41",
						   32999 => x"4c",
						   33000 => x"3f",
						   33001 => x"00",
						   33002 => x"40",
						   33003 => x"ff",
						   33004 => x"62",
						   33005 => x"51",
						   33006 => x"4f",
						   33007 => x"50",
						   33008 => x"61",
						   33009 => x"60",
						   33010 => x"70",
						   33011 => x"00",
						   33012 => x"17",
						   33013 => x"01",
						   33014 => x"00",
						   33015 => x"3d",
						   33016 => x"0a",
						   33017 => x"e2",
						   33018 => x"01",
						   33019 => x"0f",
						   33020 => x"40",
						   33021 => x"ff",
						   33022 => x"f0",
						   33023 => x"00",
						   33024 => x"ac",
						   33025 => x"81",
						   33026 => x"78",
						   33027 => x"83",
						   33028 => x"00",
						   33029 => x"80",
						   33030 => x"00",
						   33031 => x"20",
						   -- Begin: program memory TEXT Section
						   33032 => x"21",		-- 008108: 2183             DECD.W  SP
						   33033 => x"A3",
						   33034 => x"B2",		-- 00810a: B240             MOV.W   #0x5a80,&WDTCTL_L
						   33035 => x"60",
						   33036 => x"80",		-- 00810c: 805A            
						   33037 => x"5A",
						   33038 => x"CC",		-- 00810e: CC01            
						   33039 => x"01",
						   33040 => x"92",		-- 008110: 92C3             BIC.W   #1,&PM5CTL0_L
						   33041 => x"E3",
						   33042 => x"30",		-- 008112: 3001            
						   33043 => x"01",
						   33044 => x"5F",		-- 008114: 5F42             MOV.B   &P1DIR,R15
						   33045 => x"62",
						   33046 => x"04",		-- 008116: 0402            
						   33047 => x"02",
						   33048 => x"C2",		-- 008118: C243             CLR.B   &P1DIR
						   33049 => x"63",
						   33050 => x"04",		-- 00811a: 0402            
						   33051 => x"02",
						   33052 => x"F2",		-- 00811c: F2F0             AND.B   #0x00fc,&P2DIR
						   33053 => x"10",
						   33054 => x"FC",		-- 00811e: FC00            
						   33055 => x"00",
						   33056 => x"05",		-- 008120: 0502            
						   33057 => x"02",
						   33058 => x"F2",		-- 008122: F2D0             BIS.B   #0x0034,&P2DIR
						   33059 => x"F0",
						   33060 => x"34",		-- 008124: 3400            
						   33061 => x"00",
						   33062 => x"05",		-- 008126: 0502            
						   33063 => x"02",
						   33064 => x"3F",		-- 008128: 3F40             MOV.W   #0x0003,R15
						   33065 => x"60",
						   33066 => x"03",		-- 00812a: 0300            
						   33067 => x"00",
						   33068 => x"5F",		-- 00812c: 5FF2             AND.B   &P2IN,R15
						   33069 => x"12",
						   33070 => x"01",		-- 00812e: 0102            
						   33071 => x"02",
						   33072 => x"C1",		-- 008130: C14F             MOV.B   R15,0x0000(SP)
						   33073 => x"6F",
						   33074 => x"00",		-- 008132: 0000            
						   33075 => x"00",
						   33076 => x"D1",		-- 008134: D193             CMP.B   #1,0x0000(SP)
						   33077 => x"B3",
						   33078 => x"00",		-- 008136: 0000            
						   33079 => x"00",
						   33080 => x"04",		-- 008138: 0420             JNE     ($C$L8)
						   33081 => x"40",
						   33082 => x"B2",		-- 00813a: B240             MOV.W   #0x002f,&set_angle
						   33083 => x"60",
						   33084 => x"2F",		-- 00813c: 2F00            
						   33085 => x"00",
						   33086 => x"02",		-- 00813e: 0221            
						   33087 => x"21",
						   33088 => x"0A",		-- 008140: 0A3C             JMP     ($C$L10)
						   33089 => x"5C",
						   33090 => x"E1",		-- 008142: E193             CMP.B   #2,0x0000(SP)
						   33091 => x"B3",
						   33092 => x"00",		-- 008144: 0000            
						   33093 => x"00",
						   33094 => x"04",		-- 008146: 0420             JNE     ($C$L9)
						   33095 => x"40",
						   33096 => x"B2",		-- 008148: B240             MOV.W   #0x004f,&set_angle
						   33097 => x"60",
						   33098 => x"4F",		-- 00814a: 4F00            
						   33099 => x"00",
						   33100 => x"02",		-- 00814c: 0221            
						   33101 => x"21",
						   33102 => x"03",		-- 00814e: 033C             JMP     ($C$L10)
						   33103 => x"5C",
						   33104 => x"B2",		-- 008150: B240             MOV.W   #0x003d,&set_angle
						   33105 => x"60",
						   33106 => x"3D",		-- 008152: 3D00            
						   33107 => x"00",
						   33108 => x"02",		-- 008154: 0221            
						   33109 => x"21",
						   33110 => x"5F",		-- 008156: 5F42             MOV.B   &P1IN,R15
						   33111 => x"62",
						   33112 => x"00",		-- 008158: 0002            
						   33113 => x"02",
						   33114 => x"D1",		-- 00815a: D14F             MOV.B   0x2000(R15),0x0000(SP)
						   33115 => x"6F",
						   33116 => x"00",		-- 00815c: 0020            
						   33117 => x"20",
						   33118 => x"00",		-- 00815e: 0000            
						   33119 => x"00",
						   33120 => x"6F",		-- 008160: 6F41             MOV.B   @SP,R15
						   33121 => x"61",
						   33122 => x"1F",		-- 008162: 1F92             CMP.W   &set_angle,R15
						   33123 => x"B2",
						   33124 => x"02",		-- 008164: 0221            
						   33125 => x"21",
						   33126 => x"0B",		-- 008166: 0B2C             JHS     ($C$L11)
						   33127 => x"4C",
						   33128 => x"E2",		-- 008168: E2C2             BIC.B   #4,&P2OUT
						   33129 => x"E2",
						   33130 => x"03",		-- 00816a: 0302            
						   33131 => x"02",
						   33132 => x"F2",		-- 00816c: F2F0             AND.B   #0x00df,&P2OUT
						   33133 => x"10",
						   33134 => x"DF",		-- 00816e: DF00            
						   33135 => x"00",
						   33136 => x"03",		-- 008170: 0302            
						   33137 => x"02",
						   33138 => x"5F",		-- 008172: 5F42             MOV.B   &set_angle,R15
						   33139 => x"62",
						   33140 => x"02",		-- 008174: 0221            
						   33141 => x"21",
						   33142 => x"6F",		-- 008176: 6F81             SUB.B   @SP,R15
						   33143 => x"A1",
						   33144 => x"C1",		-- 008178: C14F             MOV.B   R15,0x0000(SP)
						   33145 => x"6F",
						   33146 => x"00",		-- 00817a: 0000            
						   33147 => x"00",
						   33148 => x"11",		-- 00817c: 113C             JMP     ($C$L13)
						   33149 => x"5C",
						   33150 => x"6F",		-- 00817e: 6F41             MOV.B   @SP,R15
						   33151 => x"61",
						   33152 => x"82",		-- 008180: 829F             CMP.W   R15,&set_angle
						   33153 => x"BF",
						   33154 => x"02",		-- 008182: 0221            
						   33155 => x"21",
						   33156 => x"09",		-- 008184: 092C             JHS     ($C$L12)
						   33157 => x"4C",
						   33158 => x"E2",		-- 008186: E2C2             BIC.B   #4,&P2OUT
						   33159 => x"E2",
						   33160 => x"03",		-- 008188: 0302            
						   33161 => x"02",
						   33162 => x"F2",		-- 00818a: F2D0             BIS.B   #0x0020,&P2OUT
						   33163 => x"F0",
						   33164 => x"20",		-- 00818c: 2000            
						   33165 => x"00",
						   33166 => x"03",		-- 00818e: 0302            
						   33167 => x"02",
						   33168 => x"D1",		-- 008190: D182             SUB.B   &set_angle,0x0000(SP)
						   33169 => x"A2",
						   33170 => x"02",		-- 008192: 0221            
						   33171 => x"21",
						   33172 => x"00",		-- 008194: 0000            
						   33173 => x"00",
						   33174 => x"04",		-- 008196: 043C             JMP     ($C$L13)
						   33175 => x"5C",
						   33176 => x"E2",		-- 008198: E2D2             BIS.B   #4,&P2OUT
						   33177 => x"F2",
						   33178 => x"03",		-- 00819a: 0302            
						   33179 => x"02",
						   33180 => x"C1",		-- 00819c: C143             CLR.B   0x0000(SP)
						   33181 => x"63",
						   33182 => x"00",		-- 00819e: 0000            
						   33183 => x"00",
						   33184 => x"6F",		-- 0081a0: 6F41             MOV.B   @SP,R15
						   33185 => x"61",
						   33186 => x"82",		-- 0081a2: 824F             MOV.W   R15,&frequency
						   33187 => x"6F",
						   33188 => x"00",		-- 0081a4: 0021            
						   33189 => x"21",
						   33190 => x"B0",		-- 0081a6: B012             CALL    #delay
						   33191 => x"32",
						   33192 => x"28",		-- 0081a8: 2882            
						   33193 => x"82",
						   33194 => x"BE",		-- 0081aa: BE3F             JMP     ($C$L7)
						   33195 => x"5F",
						   -- Begin: __TI_decompress_lzss
						   33196 => x"0A",		-- 0081ac: 0A12             PUSH    R10
						   33197 => x"32",
						   33198 => x"09",		-- 0081ae: 0912             PUSH    R9
						   33199 => x"32",
						   33200 => x"08",		-- 0081b0: 0812             PUSH    R8
						   33201 => x"32",
						   33202 => x"0A",		-- 0081b2: 0A4C             MOV.W   R12,R10
						   33203 => x"6C",
						   33204 => x"78",		-- 0081b4: 784A             MOV.B   @R10+,R8
						   33205 => x"6A",
						   33206 => x"09",		-- 0081b6: 0943             CLR.W   R9
						   33207 => x"63",
						   33208 => x"11",		-- 0081b8: 113C             JMP     ($C$L6)
						   33209 => x"5C",
						   33210 => x"0E",		-- 0081ba: 0E4D             MOV.W   R13,R14
						   33211 => x"6D",
						   33212 => x"0E",		-- 0081bc: 0E8B             SUB.W   R11,R14
						   33213 => x"AB",
						   33214 => x"1E",		-- 0081be: 1E83             DEC.W   R14
						   33215 => x"A3",
						   33216 => x"1D",		-- 0081c0: 1D53             INC.W   R13
						   33217 => x"73",
						   33218 => x"FD",		-- 0081c2: FD4E             MOV.B   @R14+,0xffff(R13)
						   33219 => x"6E",
						   33220 => x"FF",		-- 0081c4: FFFF            
						   33221 => x"FF",
						   33222 => x"1F",		-- 0081c6: 1F83             DEC.W   R15
						   33223 => x"A3",
						   33224 => x"FB",		-- 0081c8: FB23             JNE     ($C$L3)
						   33225 => x"43",
						   33226 => x"03",		-- 0081ca: 033C             JMP     ($C$L5)
						   33227 => x"5C",
						   33228 => x"1D",		-- 0081cc: 1D53             INC.W   R13
						   33229 => x"73",
						   33230 => x"FD",		-- 0081ce: FD4A             MOV.B   @R10+,0xffff(R13)
						   33231 => x"6A",
						   33232 => x"FF",		-- 0081d0: FFFF            
						   33233 => x"FF",
						   33234 => x"12",		-- 0081d2: 12C3             CLRC    
						   33235 => x"E3",
						   33236 => x"08",		-- 0081d4: 0810             RRC     R8
						   33237 => x"30",
						   33238 => x"19",		-- 0081d6: 1953             INC.W   R9
						   33239 => x"73",
						   33240 => x"39",		-- 0081d8: 3992             CMP.W   #8,R9
						   33241 => x"B2",
						   33242 => x"EC",		-- 0081da: EC37             JGE     ($C$L1)
						   33243 => x"57",
						   33244 => x"18",		-- 0081dc: 18B3             BIT.W   #1,R8
						   33245 => x"D3",
						   33246 => x"F6",		-- 0081de: F623             JNE     ($C$L4)
						   33247 => x"43",
						   33248 => x"7B",		-- 0081e0: 7B4A             MOV.B   @R10+,R11
						   33249 => x"6A",
						   33250 => x"7F",		-- 0081e2: 7F4A             MOV.B   @R10+,R15
						   33251 => x"6A",
						   33252 => x"0C",		-- 0081e4: 0C4B             MOV.W   R11,R12
						   33253 => x"6B",
						   33254 => x"B0",		-- 0081e6: B012             CALL    #__mspabi_slli_4
						   33255 => x"32",
						   33256 => x"52",		-- 0081e8: 5283            
						   33257 => x"83",
						   33258 => x"0B",		-- 0081ea: 0B4C             MOV.W   R12,R11
						   33259 => x"6C",
						   33260 => x"0C",		-- 0081ec: 0C4F             MOV.W   R15,R12
						   33261 => x"6F",
						   33262 => x"B0",		-- 0081ee: B012             CALL    #__mspabi_srli_4
						   33263 => x"32",
						   33264 => x"DC",		-- 0081f0: DC82            
						   33265 => x"82",
						   33266 => x"3C",		-- 0081f2: 3CF0             AND.W   #0x000f,R12
						   33267 => x"10",
						   33268 => x"0F",		-- 0081f4: 0F00            
						   33269 => x"00",
						   33270 => x"0B",		-- 0081f6: 0BDC             BIS.W   R12,R11
						   33271 => x"FC",
						   33272 => x"3F",		-- 0081f8: 3FF0             AND.W   #0x000f,R15
						   33273 => x"10",
						   33274 => x"0F",		-- 0081fa: 0F00            
						   33275 => x"00",
						   33276 => x"3F",		-- 0081fc: 3F50             ADD.W   #0x0003,R15
						   33277 => x"70",
						   33278 => x"03",		-- 0081fe: 0300            
						   33279 => x"00",
						   33280 => x"3F",		-- 008200: 3F90             CMP.W   #0x0012,R15
						   33281 => x"B0",
						   33282 => x"12",		-- 008202: 1200            
						   33283 => x"00",
						   33284 => x"0C",		-- 008204: 0C20             JNE     ($C$L8)
						   33285 => x"40",
						   33286 => x"7E",		-- 008206: 7E4A             MOV.B   @R10+,R14
						   33287 => x"6A",
						   33288 => x"3E",		-- 008208: 3EB0             BIT.W   #0x0080,R14
						   33289 => x"D0",
						   33290 => x"80",		-- 00820a: 8000            
						   33291 => x"00",
						   33292 => x"07",		-- 00820c: 0724             JEQ     ($C$L7)
						   33293 => x"44",
						   33294 => x"7C",		-- 00820e: 7C4A             MOV.B   @R10+,R12
						   33295 => x"6A",
						   33296 => x"4C",		-- 008210: 4C4C             MOV.B   R12,R12
						   33297 => x"6C",
						   33298 => x"B0",		-- 008212: B012             CALL    #__mspabi_slli_7
						   33299 => x"32",
						   33300 => x"4C",		-- 008214: 4C83            
						   33301 => x"83",
						   33302 => x"3E",		-- 008216: 3EF0             AND.W   #0x007f,R14
						   33303 => x"10",
						   33304 => x"7F",		-- 008218: 7F00            
						   33305 => x"00",
						   33306 => x"0E",		-- 00821a: 0EDC             BIS.W   R12,R14
						   33307 => x"FC",
						   33308 => x"0F",		-- 00821c: 0F5E             ADD.W   R14,R15
						   33309 => x"7E",
						   33310 => x"3B",		-- 00821e: 3B90             CMP.W   #0x0fff,R11
						   33311 => x"B0",
						   33312 => x"FF",		-- 008220: FF0F            
						   33313 => x"0F",
						   33314 => x"CB",		-- 008222: CB23             JNE     ($C$L2)
						   33315 => x"43",
						   33316 => x"30",		-- 008224: 3040             BR      #__mspabi_func_epilog_3
						   33317 => x"60",
						   33318 => x"A4",		-- 008226: A483            
						   33319 => x"83",
						   -- Begin: delay
						   33320 => x"92",		-- 008228: 9253             INC.W   &delayCounter
						   33321 => x"73",
						   33322 => x"04",		-- 00822a: 0421            
						   33323 => x"21",
						   33324 => x"82",		-- 00822c: 8263             ADC.W   &0x2106
						   33325 => x"83",
						   33326 => x"06",		-- 00822e: 0621            
						   33327 => x"21",
						   33328 => x"92",		-- 008230: 9292             CMP.W   &0x210a,&0x2106
						   33329 => x"B2",
						   33330 => x"0A",		-- 008232: 0A21            
						   33331 => x"21",
						   33332 => x"06",		-- 008234: 0621            
						   33333 => x"21",
						   33334 => x"34",		-- 008236: 3428             JLO     ($C$L6)
						   33335 => x"48",
						   33336 => x"04",		-- 008238: 0420             JNE     ($C$L1)
						   33337 => x"40",
						   33338 => x"92",		-- 00823a: 9292             CMP.W   &delayLength,&delayCounter
						   33339 => x"B2",
						   33340 => x"08",		-- 00823c: 0821            
						   33341 => x"21",
						   33342 => x"04",		-- 00823e: 0421            
						   33343 => x"21",
						   33344 => x"2F",		-- 008240: 2F28             JLO     ($C$L6)
						   33345 => x"48",
						   33346 => x"82",		-- 008242: 8293             TST.W   &frequency
						   33347 => x"B3",
						   33348 => x"00",		-- 008244: 0021            
						   33349 => x"21",
						   33350 => x"04",		-- 008246: 0434             JGE     ($C$L2)
						   33351 => x"54",
						   33352 => x"B2",		-- 008248: B2E3             INV.W   &frequency
						   33353 => x"03",
						   33354 => x"00",		-- 00824a: 0021            
						   33355 => x"21",
						   33356 => x"92",		-- 00824c: 9253             INC.W   &frequency
						   33357 => x"73",
						   33358 => x"00",		-- 00824e: 0021            
						   33359 => x"21",
						   33360 => x"1E",		-- 008250: 1E42             MOV.W   &frequency,R14
						   33361 => x"62",
						   33362 => x"00",		-- 008252: 0021            
						   33363 => x"21",
						   33364 => x"3E",		-- 008254: 3EB0             BIT.W   #0x8000,R14
						   33365 => x"D0",
						   33366 => x"00",		-- 008256: 0080            
						   33367 => x"80",
						   33368 => x"0F",		-- 008258: 0F7F             SUBC.W  R15,R15
						   33369 => x"9F",
						   33370 => x"3F",		-- 00825a: 3FE3             INV.W   R15
						   33371 => x"03",
						   33372 => x"82",		-- 00825c: 824E             MOV.W   R14,&delayLength
						   33373 => x"6E",
						   33374 => x"08",		-- 00825e: 0821            
						   33375 => x"21",
						   33376 => x"82",		-- 008260: 824F             MOV.W   R15,&0x210a
						   33377 => x"6F",
						   33378 => x"0A",		-- 008262: 0A21            
						   33379 => x"21",
						   33380 => x"82",		-- 008264: 8293             TST.W   &0x210a
						   33381 => x"B3",
						   33382 => x"0A",		-- 008266: 0A21            
						   33383 => x"21",
						   33384 => x"04",		-- 008268: 0420             JNE     ($C$L3)
						   33385 => x"40",
						   33386 => x"B2",		-- 00826a: B290             CMP.W   #0x000e,&delayLength
						   33387 => x"B0",
						   33388 => x"0E",		-- 00826c: 0E00            
						   33389 => x"00",
						   33390 => x"08",		-- 00826e: 0821            
						   33391 => x"21",
						   33392 => x"06",		-- 008270: 0628             JLO     ($C$L4)
						   33393 => x"48",
						   33394 => x"B2",		-- 008272: B240             MOV.W   #0x000d,&delayLength
						   33395 => x"60",
						   33396 => x"0D",		-- 008274: 0D00            
						   33397 => x"00",
						   33398 => x"08",		-- 008276: 0821            
						   33399 => x"21",
						   33400 => x"82",		-- 008278: 8243             CLR.W   &0x210a
						   33401 => x"63",
						   33402 => x"0A",		-- 00827a: 0A21            
						   33403 => x"21",
						   33404 => x"0A",		-- 00827c: 0A3C             JMP     ($C$L5)
						   33405 => x"5C",
						   33406 => x"82",		-- 00827e: 8293             TST.W   &0x210a
						   33407 => x"B3",
						   33408 => x"0A",		-- 008280: 0A21            
						   33409 => x"21",
						   33410 => x"07",		-- 008282: 0720             JNE     ($C$L5)
						   33411 => x"40",
						   33412 => x"82",		-- 008284: 8293             TST.W   &delayLength
						   33413 => x"B3",
						   33414 => x"08",		-- 008286: 0821            
						   33415 => x"21",
						   33416 => x"04",		-- 008288: 0420             JNE     ($C$L5)
						   33417 => x"40",
						   33418 => x"92",		-- 00828a: 9243             MOV.W   #1,&delayLength
						   33419 => x"63",
						   33420 => x"08",		-- 00828c: 0821            
						   33421 => x"21",
						   33422 => x"82",		-- 00828e: 8243             CLR.W   &0x210a
						   33423 => x"63",
						   33424 => x"0A",		-- 008290: 0A21            
						   33425 => x"21",
						   33426 => x"F2",		-- 008292: F2E0             XOR.B   #0x0010,&P2OUT
						   33427 => x"00",
						   33428 => x"10",		-- 008294: 1000            
						   33429 => x"00",
						   33430 => x"03",		-- 008296: 0302            
						   33431 => x"02",
						   33432 => x"82",		-- 008298: 8243             CLR.W   &delayCounter
						   33433 => x"63",
						   33434 => x"04",		-- 00829a: 0421            
						   33435 => x"21",
						   33436 => x"82",		-- 00829c: 8243             CLR.W   &0x2106
						   33437 => x"63",
						   33438 => x"06",		-- 00829e: 0621            
						   33439 => x"21",
						   33440 => x"30",		-- 0082a0: 3041             RET     
						   33441 => x"61",
						   -- Begin: __mspabi_srli
						   33442 => x"3D",		-- 0082a2: 3DF0             AND.W   #0x000f,R13
						   33443 => x"10",
						   33444 => x"0F",		-- 0082a4: 0F00            
						   33445 => x"00",
						   33446 => x"3D",		-- 0082a6: 3DE0             XOR.W   #0x000f,R13
						   33447 => x"00",
						   33448 => x"0F",		-- 0082a8: 0F00            
						   33449 => x"00",
						   33450 => x"0D",		-- 0082aa: 0D5D             RLA.W   R13
						   33451 => x"7D",
						   33452 => x"0D",		-- 0082ac: 0D5D             RLA.W   R13
						   33453 => x"7D",
						   33454 => x"00",		-- 0082ae: 005D             ADD.W   R13,PC
						   33455 => x"7D",
						   -- Begin: __mspabi_srli_15
						   33456 => x"12",		-- 0082b0: 12C3             CLRC    
						   33457 => x"E3",
						   33458 => x"0C",		-- 0082b2: 0C10             RRC     R12
						   33459 => x"30",
						   -- Begin: __mspabi_srli_14
						   33460 => x"12",		-- 0082b4: 12C3             CLRC    
						   33461 => x"E3",
						   33462 => x"0C",		-- 0082b6: 0C10             RRC     R12
						   33463 => x"30",
						   -- Begin: __mspabi_srli_13
						   33464 => x"12",		-- 0082b8: 12C3             CLRC    
						   33465 => x"E3",
						   33466 => x"0C",		-- 0082ba: 0C10             RRC     R12
						   33467 => x"30",
						   -- Begin: __mspabi_srli_12
						   33468 => x"12",		-- 0082bc: 12C3             CLRC    
						   33469 => x"E3",
						   33470 => x"0C",		-- 0082be: 0C10             RRC     R12
						   33471 => x"30",
						   -- Begin: __mspabi_srli_11
						   33472 => x"12",		-- 0082c0: 12C3             CLRC    
						   33473 => x"E3",
						   33474 => x"0C",		-- 0082c2: 0C10             RRC     R12
						   33475 => x"30",
						   -- Begin: __mspabi_srli_10
						   33476 => x"12",		-- 0082c4: 12C3             CLRC    
						   33477 => x"E3",
						   33478 => x"0C",		-- 0082c6: 0C10             RRC     R12
						   33479 => x"30",
						   -- Begin: __mspabi_srli_9
						   33480 => x"12",		-- 0082c8: 12C3             CLRC    
						   33481 => x"E3",
						   33482 => x"0C",		-- 0082ca: 0C10             RRC     R12
						   33483 => x"30",
						   -- Begin: __mspabi_srli_8
						   33484 => x"12",		-- 0082cc: 12C3             CLRC    
						   33485 => x"E3",
						   33486 => x"0C",		-- 0082ce: 0C10             RRC     R12
						   33487 => x"30",
						   -- Begin: __mspabi_srli_7
						   33488 => x"12",		-- 0082d0: 12C3             CLRC    
						   33489 => x"E3",
						   33490 => x"0C",		-- 0082d2: 0C10             RRC     R12
						   33491 => x"30",
						   -- Begin: __mspabi_srli_6
						   33492 => x"12",		-- 0082d4: 12C3             CLRC    
						   33493 => x"E3",
						   33494 => x"0C",		-- 0082d6: 0C10             RRC     R12
						   33495 => x"30",
						   -- Begin: __mspabi_srli_5
						   33496 => x"12",		-- 0082d8: 12C3             CLRC    
						   33497 => x"E3",
						   33498 => x"0C",		-- 0082da: 0C10             RRC     R12
						   33499 => x"30",
						   -- Begin: __mspabi_srli_4
						   33500 => x"12",		-- 0082dc: 12C3             CLRC    
						   33501 => x"E3",
						   33502 => x"0C",		-- 0082de: 0C10             RRC     R12
						   33503 => x"30",
						   -- Begin: __mspabi_srli_3
						   33504 => x"12",		-- 0082e0: 12C3             CLRC    
						   33505 => x"E3",
						   33506 => x"0C",		-- 0082e2: 0C10             RRC     R12
						   33507 => x"30",
						   -- Begin: __mspabi_srli_2
						   33508 => x"12",		-- 0082e4: 12C3             CLRC    
						   33509 => x"E3",
						   33510 => x"0C",		-- 0082e6: 0C10             RRC     R12
						   33511 => x"30",
						   -- Begin: __mspabi_srli_1
						   33512 => x"12",		-- 0082e8: 12C3             CLRC    
						   33513 => x"E3",
						   33514 => x"0C",		-- 0082ea: 0C10             RRC     R12
						   33515 => x"30",
						   33516 => x"30",		-- 0082ec: 3041             RET     
						   33517 => x"61",
						   -- Begin: __TI_auto_init_nobinit_nopinit
						   33518 => x"0A",		-- 0082ee: 0A12             PUSH    R10
						   33519 => x"32",
						   33520 => x"09",		-- 0082f0: 0912             PUSH    R9
						   33521 => x"32",
						   33522 => x"3F",		-- 0082f2: 3F40             MOV.W   #0x8100,R15
						   33523 => x"60",
						   33524 => x"00",		-- 0082f4: 0081            
						   33525 => x"81",
						   33526 => x"3F",		-- 0082f6: 3F90             CMP.W   #0x8104,R15
						   33527 => x"B0",
						   33528 => x"04",		-- 0082f8: 0481            
						   33529 => x"81",
						   33530 => x"16",		-- 0082fa: 1624             JEQ     ($C$L22)
						   33531 => x"44",
						   33532 => x"3F",		-- 0082fc: 3F40             MOV.W   #0x8104,R15
						   33533 => x"60",
						   33534 => x"04",		-- 0082fe: 0481            
						   33535 => x"81",
						   33536 => x"3F",		-- 008300: 3F90             CMP.W   #0x8108,R15
						   33537 => x"B0",
						   33538 => x"08",		-- 008302: 0881            
						   33539 => x"81",
						   33540 => x"11",		-- 008304: 1124             JEQ     ($C$L22)
						   33541 => x"44",
						   33542 => x"3A",		-- 008306: 3A40             MOV.W   #0x8108,R10
						   33543 => x"60",
						   33544 => x"08",		-- 008308: 0881            
						   33545 => x"81",
						   33546 => x"3A",		-- 00830a: 3A80             SUB.W   #0x8104,R10
						   33547 => x"A0",
						   33548 => x"04",		-- 00830c: 0481            
						   33549 => x"81",
						   33550 => x"0A",		-- 00830e: 0A11             RRA     R10
						   33551 => x"31",
						   33552 => x"0A",		-- 008310: 0A11             RRA     R10
						   33553 => x"31",
						   33554 => x"39",		-- 008312: 3940             MOV.W   #0x8104,R9
						   33555 => x"60",
						   33556 => x"04",		-- 008314: 0481            
						   33557 => x"81",
						   33558 => x"3C",		-- 008316: 3C49             MOV.W   @R9+,R12
						   33559 => x"69",
						   33560 => x"7F",		-- 008318: 7F4C             MOV.B   @R12+,R15
						   33561 => x"6C",
						   33562 => x"0F",		-- 00831a: 0F5F             RLA.W   R15
						   33563 => x"7F",
						   33564 => x"1F",		-- 00831c: 1F4F             MOV.W   0x8100(R15),R15
						   33565 => x"6F",
						   33566 => x"00",		-- 00831e: 0081            
						   33567 => x"81",
						   33568 => x"3D",		-- 008320: 3D49             MOV.W   @R9+,R13
						   33569 => x"69",
						   33570 => x"8F",		-- 008322: 8F12             CALL    R15
						   33571 => x"32",
						   33572 => x"1A",		-- 008324: 1A83             DEC.W   R10
						   33573 => x"A3",
						   33574 => x"F7",		-- 008326: F723             JNE     ($C$L21)
						   33575 => x"43",
						   33576 => x"B0",		-- 008328: B012             CALL    #_system_post_cinit
						   33577 => x"32",
						   33578 => x"B6",		-- 00832a: B683            
						   33579 => x"83",
						   33580 => x"30",		-- 00832c: 3040             BR      #__mspabi_func_epilog_2
						   33581 => x"60",
						   33582 => x"A6",		-- 00832e: A683            
						   33583 => x"83",
						   -- Begin: __mspabi_slli
						   33584 => x"3D",		-- 008330: 3DF0             AND.W   #0x000f,R13
						   33585 => x"10",
						   33586 => x"0F",		-- 008332: 0F00            
						   33587 => x"00",
						   33588 => x"3D",		-- 008334: 3DE0             XOR.W   #0x000f,R13
						   33589 => x"00",
						   33590 => x"0F",		-- 008336: 0F00            
						   33591 => x"00",
						   33592 => x"0D",		-- 008338: 0D5D             RLA.W   R13
						   33593 => x"7D",
						   33594 => x"00",		-- 00833a: 005D             ADD.W   R13,PC
						   33595 => x"7D",
						   -- Begin: __mspabi_slli_15
						   33596 => x"0C",		-- 00833c: 0C5C             RLA.W   R12
						   33597 => x"7C",
						   -- Begin: __mspabi_slli_14
						   33598 => x"0C",		-- 00833e: 0C5C             RLA.W   R12
						   33599 => x"7C",
						   -- Begin: __mspabi_slli_13
						   33600 => x"0C",		-- 008340: 0C5C             RLA.W   R12
						   33601 => x"7C",
						   -- Begin: __mspabi_slli_12
						   33602 => x"0C",		-- 008342: 0C5C             RLA.W   R12
						   33603 => x"7C",
						   -- Begin: __mspabi_slli_11
						   33604 => x"0C",		-- 008344: 0C5C             RLA.W   R12
						   33605 => x"7C",
						   -- Begin: __mspabi_slli_10
						   33606 => x"0C",		-- 008346: 0C5C             RLA.W   R12
						   33607 => x"7C",
						   -- Begin: __mspabi_slli_9
						   33608 => x"0C",		-- 008348: 0C5C             RLA.W   R12
						   33609 => x"7C",
						   -- Begin: __mspabi_slli_8
						   33610 => x"0C",		-- 00834a: 0C5C             RLA.W   R12
						   33611 => x"7C",
						   -- Begin: __mspabi_slli_7
						   33612 => x"0C",		-- 00834c: 0C5C             RLA.W   R12
						   33613 => x"7C",
						   -- Begin: __mspabi_slli_6
						   33614 => x"0C",		-- 00834e: 0C5C             RLA.W   R12
						   33615 => x"7C",
						   -- Begin: __mspabi_slli_5
						   33616 => x"0C",		-- 008350: 0C5C             RLA.W   R12
						   33617 => x"7C",
						   -- Begin: __mspabi_slli_4
						   33618 => x"0C",		-- 008352: 0C5C             RLA.W   R12
						   33619 => x"7C",
						   -- Begin: __mspabi_slli_3
						   33620 => x"0C",		-- 008354: 0C5C             RLA.W   R12
						   33621 => x"7C",
						   -- Begin: __mspabi_slli_2
						   33622 => x"0C",		-- 008356: 0C5C             RLA.W   R12
						   33623 => x"7C",
						   -- Begin: __mspabi_slli_1
						   33624 => x"0C",		-- 008358: 0C5C             RLA.W   R12
						   33625 => x"7C",
						   33626 => x"30",		-- 00835a: 3041             RET     
						   33627 => x"61",
						   -- Begin: _c_int00_noargs
						   33628 => x"31",		-- 00835c: 3140             MOV.W   #0x3000,SP
						   33629 => x"60",
						   33630 => x"00",		-- 00835e: 0030            
						   33631 => x"30",
						   33632 => x"B0",		-- 008360: B012             CALL    #_system_pre_init
						   33633 => x"32",
						   33634 => x"B2",		-- 008362: B283            
						   33635 => x"83",
						   33636 => x"0C",		-- 008364: 0C93             TST.W   R12
						   33637 => x"B3",
						   33638 => x"02",		-- 008366: 0224             JEQ     ($C$L2)
						   33639 => x"44",
						   33640 => x"B0",		-- 008368: B012             CALL    #__TI_auto_init_nobinit_nopinit
						   33641 => x"32",
						   33642 => x"EE",		-- 00836a: EE82            
						   33643 => x"82",
						   33644 => x"0C",		-- 00836c: 0C43             CLR.W   R12
						   33645 => x"63",
						   33646 => x"B0",		-- 00836e: B012             CALL    #main
						   33647 => x"32",
						   33648 => x"08",		-- 008370: 0881            
						   33649 => x"81",
						   33650 => x"1C",		-- 008372: 1C43             MOV.W   #1,R12
						   33651 => x"63",
						   33652 => x"B0",		-- 008374: B012             CALL    #abort
						   33653 => x"32",
						   33654 => x"AC",		-- 008376: AC83            
						   33655 => x"83",
						   -- Begin: __TI_decompress_none
						   33656 => x"0F",		-- 008378: 0F4C             MOV.W   R12,R15
						   33657 => x"6C",
						   33658 => x"0C",		-- 00837a: 0C4D             MOV.W   R13,R12
						   33659 => x"6D",
						   33660 => x"3D",		-- 00837c: 3D40             MOV.W   #0x0003,R13
						   33661 => x"60",
						   33662 => x"03",		-- 00837e: 0300            
						   33663 => x"00",
						   33664 => x"0D",		-- 008380: 0D5F             ADD.W   R15,R13
						   33665 => x"7F",
						   33666 => x"1E",		-- 008382: 1E4F             MOV.W   0x0001(R15),R14
						   33667 => x"6F",
						   33668 => x"01",		-- 008384: 0100            
						   33669 => x"00",
						   33670 => x"30",		-- 008386: 3040             BR      #memcpy
						   33671 => x"60",
						   33672 => x"8A",		-- 008388: 8A83            
						   33673 => x"83",
						   -- Begin: memcpy
						   33674 => x"0E",		-- 00838a: 0E93             TST.W   R14
						   33675 => x"B3",
						   33676 => x"06",		-- 00838c: 0624             JEQ     ($C$L2)
						   33677 => x"44",
						   33678 => x"0F",		-- 00838e: 0F4C             MOV.W   R12,R15
						   33679 => x"6C",
						   33680 => x"1F",		-- 008390: 1F53             INC.W   R15
						   33681 => x"73",
						   33682 => x"FF",		-- 008392: FF4D             MOV.B   @R13+,0xffff(R15)
						   33683 => x"6D",
						   33684 => x"FF",		-- 008394: FFFF            
						   33685 => x"FF",
						   33686 => x"1E",		-- 008396: 1E83             DEC.W   R14
						   33687 => x"A3",
						   33688 => x"FB",		-- 008398: FB23             JNE     ($C$L1)
						   33689 => x"43",
						   33690 => x"30",		-- 00839a: 3041             RET     
						   33691 => x"61",
						   -- Begin: __mspabi_func_epilog_7
						   -- Begin: __mspabi_func_epilog
						   33692 => x"34",		-- 00839c: 3441             POP.W   R4
						   33693 => x"61",
						   -- Begin: __mspabi_func_epilog_6
						   33694 => x"35",		-- 00839e: 3541             POP.W   R5
						   33695 => x"61",
						   -- Begin: __mspabi_func_epilog_5
						   33696 => x"36",		-- 0083a0: 3641             POP.W   R6
						   33697 => x"61",
						   -- Begin: __mspabi_func_epilog_4
						   33698 => x"37",		-- 0083a2: 3741             POP.W   R7
						   33699 => x"61",
						   -- Begin: __mspabi_func_epilog_3
						   33700 => x"38",		-- 0083a4: 3841             POP.W   R8
						   33701 => x"61",
						   -- Begin: __mspabi_func_epilog_2
						   33702 => x"39",		-- 0083a6: 3941             POP.W   R9
						   33703 => x"61",
						   -- Begin: __mspabi_func_epilog_1
						   33704 => x"3A",		-- 0083a8: 3A41             POP.W   R10
						   33705 => x"61",
						   33706 => x"30",		-- 0083aa: 3041             RET     
						   33707 => x"61",
						   -- Begin: abort
						   33708 => x"03",		-- 0083ac: 0343             NOP     
						   33709 => x"63",
						   33710 => x"FF",		-- 0083ae: FF3F             JMP     ($C$L1)
						   33711 => x"5F",
						   33712 => x"03",		-- 0083b0: 0343             NOP     
						   33713 => x"63",
						   -- Begin: _system_pre_init
						   33714 => x"1C",		-- 0083b2: 1C43             MOV.W   #1,R12
						   33715 => x"63",
						   33716 => x"30",		-- 0083b4: 3041             RET     
						   33717 => x"61",
						   -- Begin: _system_post_cinit
						   33718 => x"30",		-- 0083b6: 3041             RET     
						   33719 => x"61",
						   -- ISR Trap
						   33720 => x"32",		-- 0083b8: 32D0             BIS.W   #0x0010,SR
						   33721 => x"F0",
						   33722 => x"10",		-- 0083ba: 1000            
						   33723 => x"00",
						   33724 => x"FD",		-- 0083bc: FD3F             JMP     (__TI_ISR_TRAP)
						   33725 => x"5F",
						   33726 => x"03",		-- 0083be: 0343             NOP     
						   33727 => x"63",
						   -- IRQ Vectors (Interrupt Vectors)
						   65486 => x"b8",		-- 00ffce:83b8 PORT4 __TI_int22 int22
						   65487 => x"83",
						   65488 => x"b8",		-- 00ffd0:83b8 PORT3 __TI_int23 int23
						   65489 => x"83",
						   65490 => x"b8",		-- 00ffd2:83b8 PORT2 __TI_int24 int24
						   65491 => x"83",
						   65492 => x"b8",		-- 00ffd4:83b8 PORT1 __TI_int25 int25
						   65493 => x"83",
						   65494 => x"b8",		-- 00ffd6:83b8 SAC1_SAC3 __TI_int26 int26
						   65495 => x"83",
						   65496 => x"b8",		-- 00ffd8:83b8 SAC0_SAC2 __TI_int27 int27
						   65497 => x"83",
						   65498 => x"b8",		-- 00ffda:83b8 ECOMP0_ECOMP1 __TI_int28 int28
						   65499 => x"83",
						   65500 => x"b8",		-- 00ffdc:83b8 ADC __TI_int29 int29
						   65501 => x"83",
						   65502 => x"b8",		-- 00ffde:83b8 EUSCI_B1 __TI_int30 int30
						   65503 => x"83",
						   65504 => x"b8",		-- 00ffe0:83b8 EUSCI_B0 __TI_int31 int31
						   65505 => x"83",
						   65506 => x"b8",		-- 00ffe2:83b8 EUSCI_A1 __TI_int32 int32
						   65507 => x"83",
						   65508 => x"b8",		-- 00ffe4:83b8 EUSCI_A0 __TI_int33 int33
						   65509 => x"83",
						   65510 => x"b8",		-- 00ffe6:83b8 WDT __TI_int34 int34
						   65511 => x"83",
						   65512 => x"b8",		-- 00ffe8:83b8 RTC __TI_int35 int35
						   65513 => x"83",
						   65514 => x"b8",		-- 00ffea:83b8 TIMER3_B1 __TI_int36 int36
						   65515 => x"83",
						   65516 => x"b8",		-- 00ffec:83b8 TIMER3_B0 __TI_int37 int37
						   65517 => x"83",
						   65518 => x"b8",		-- 00ffee:83b8 TIMER2_B1 __TI_int38 int38
						   65519 => x"83",
						   65520 => x"b8",		-- 00fff0:83b8 TIMER2_B0 __TI_int39 int39
						   65521 => x"83",
						   65522 => x"b8",		-- 00fff2:83b8 TIMER1_B1 __TI_int40 int40
						   65523 => x"83",
						   65524 => x"b8",		-- 00fff4:83b8 TIMER1_B0 __TI_int41 int41
						   65525 => x"83",
						   65526 => x"b8",		-- 00fff6:83b8 TIMER0_B1 __TI_int42 int42
						   65527 => x"83",
						   65528 => x"b8",		-- 00fff8:83b8 TIMER0_B0 __TI_int43 int43
						   65529 => x"83",
						   65530 => x"b8",		-- 00fffa:83b8 UNMI __TI_int44 int44
						   65531 => x"83",
						   65532 => x"b8",		-- 00fffc:83b8 SYSNMI __TI_int45 int45
						   65533 => x"83",
						   65534 => x"5c",		-- 00fffe:835c .reset _reset_vector reset
						   65535 => x"83",
						   others => x"00");

    signal EN : std_logic;
    
    begin
    -- Note 1:  The bus system uses a 16-bit Address (MAB)
    --          This address size can access locations from x0000 to xFFFF
    --          But our array is only defined from x8000 to xFFFF and
    --          if we try to access it with any other address, it will crash.
    --          So the first thing we need to do is create a local enable that
    --          will only assert when MAB is within x8000 to xFFFF.

     LOCAL_EN : process (MAB) 
     begin
         if ( (to_integer(unsigned(MAB)) >= 32768) and (to_integer(unsigned(MAB)) <= 65535)) then
           EN <= '1';
         else 
           EN <= '0';
         end if;
     end process;

    
    -- Note 2:  The bus system uses a 16-bit Address (MAB)
    --          The MDB_out is also provided as a 16-bit word
    --          However, the memory array is actually built as 8-bit bytes.
    --          So for a given 16-bit MAB, we give MDB_out = HB : LB
    --                                                 or  = ROM(MAB);1) : ROM(MAB)

    MEMORY_ROM : process (clk) 
    begin
        if (rising_edge(clk)) then
            if (EN='1' and write='0') then
                if(Byte = '0') then                      
                    MDB_in <= ROM(to_integer(unsigned(MAB)) + 1 ) & ROM(to_integer(unsigned(MAB)));
                else
                    MDB_in <= x"00" & ROM(to_integer(unsigned(MAB)));
                end if;
            end if;
        end if;
    end process;


end architecture;