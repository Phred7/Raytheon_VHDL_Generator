library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;


entity lowlife_memory is
    port ( clk	: in	std_logic;
         MAB		: in	std_logic_vector(15 downto 0);
         MDB_in  	: out	std_logic_vector(15 downto 0);
         MDB_out  	: in	std_logic_vector(15 downto 0);
         write	    : in	std_logic);
end entity;

architecture lowlife_memory_arch of lowlife_memory is

type rom_type is array (32768 to 65535) of std_logic_vector(7 downto 0);  -- this is MAB: x8000 to xFFFF
    
constant ROM : rom_type :=(						   55360 => x"B2",		-- 00d840: B240             MOV.W   #0x5a80,&WDTCTL_L
						   55361 => x"20",
						   55362 => x"80",		-- 00d842: 805A            
						   55363 => x"5A",
						   55364 => x"CC",		-- 00d844: CC01            
						   55365 => x"01",
						   55366 => x"91",		-- 00d846: 9142             MOV.W   &$P$T0$1,0x0002(SP)
						   55367 => x"22",
						   55368 => x"56",		-- 00d848: 569A            
						   55369 => x"9A",
						   55370 => x"02",		-- 00d84a: 0200            
						   55371 => x"00",
						   55372 => x"91",		-- 00d84c: 9142             MOV.W   &0x9a58,0x0004(SP)
						   55373 => x"22",
						   55374 => x"58",		-- 00d84e: 589A            
						   55375 => x"9A",
						   55376 => x"04",		-- 00d850: 0400            
						   55377 => x"00",
						   55378 => x"91",		-- 00d852: 9142             MOV.W   &0x9a5a,0x0006(SP)
						   55379 => x"22",
						   55380 => x"5A",		-- 00d854: 5A9A            
						   55381 => x"9A",
						   55382 => x"06",		-- 00d856: 0600            
						   55383 => x"00",
						   55384 => x"91",		-- 00d858: 9142             MOV.W   &0x9a5c,0x0008(SP)
						   55385 => x"22",
						   55386 => x"5C",		-- 00d85a: 5C9A            
						   55387 => x"9A",
						   55388 => x"08",		-- 00d85c: 0800            
						   55389 => x"00",
						   55390 => x"81",		-- 00d85e: 8143             CLR.W   0x000c(SP)
						   55391 => x"23",
						   55392 => x"0C",		-- 00d860: 0C00            
						   55393 => x"00",
						   55394 => x"1C",		-- 00d862: 1C41             MOV.W   0x000a(SP),R12
						   55395 => x"21",
						   55396 => x"0A",		-- 00d864: 0A00            
						   55397 => x"00",
						   55398 => x"B0",		-- 00d866: B012             CALL    #buff_value
						   55399 => x"F2",
						   55400 => x"4C",		-- 00d868: 4CE1            
						   55401 => x"E1",
						   55402 => x"1C",		-- 00d86a: 1C41             MOV.W   0x000e(SP),R12
						   55403 => x"21",
						   55404 => x"0E",		-- 00d86c: 0E00            
						   55405 => x"00",
						   55406 => x"B0",		-- 00d86e: B012             CALL    #buff_value
						   55407 => x"F2",
						   55408 => x"4C",		-- 00d870: 4CE1            
						   55409 => x"E1",
						   55410 => x"81",		-- 00d872: 8193             TST.W   0x000c(SP)
						   55411 => x"73",
						   55412 => x"0C",		-- 00d874: 0C00            
						   55413 => x"00",
						   55414 => x"06",		-- 00d876: 0620             JNE     ($C$L1)
						   55415 => x"00",
						   55416 => x"B1",		-- 00d878: B140             MOV.W   #0x852c,0x0000(SP)
						   55417 => x"20",
						   55418 => x"2C",		-- 00d87a: 2C85            
						   55419 => x"85",
						   55420 => x"00",		-- 00d87c: 0000            
						   55421 => x"00",
						   55422 => x"B0",		-- 00d87e: B012             CALL    #printf
						   55423 => x"F2",
						   55424 => x"16",		-- 00d880: 16DD            
						   55425 => x"DD",
						   55426 => x"05",		-- 00d882: 053C             JMP     ($C$L2)
						   55427 => x"1C",
						   55428 => x"B1",		-- 00d884: B140             MOV.W   #0x852c,0x0000(SP)
						   55429 => x"20",
						   55430 => x"2C",		-- 00d886: 2C85            
						   55431 => x"85",
						   55432 => x"00",		-- 00d888: 0000            
						   55433 => x"00",
						   55434 => x"B0",		-- 00d88a: B012             CALL    #printf
						   55435 => x"F2",
						   55436 => x"16",		-- 00d88c: 16DD            
						   55437 => x"DD",
						   55438 => x"0C",		-- 00d88e: 0C43             CLR.W   R12
						   55439 => x"23",
						   55440 => x"31",		-- 00d890: 3150             ADD.W   #0x0010,SP
						   55441 => x"30",
						   55442 => x"10",		-- 00d892: 1000            
						   55443 => x"00",
						   55444 => x"30",		-- 00d894: 3041             RET     
						   55445 => x"21",
						   -- Begin: getdevice
						   55446 => x"0A",		-- 00d896: 0A12             PUSH    R10
						   55447 => x"F2",
						   55448 => x"09",		-- 00d898: 0912             PUSH    R9
						   55449 => x"F2",
						   55450 => x"08",		-- 00d89a: 0812             PUSH    R8
						   55451 => x"F2",
						   55452 => x"31",		-- 00d89c: 3180             SUB.W   #0x000a,SP
						   55453 => x"60",
						   55454 => x"0A",		-- 00d89e: 0A00            
						   55455 => x"00",
						   55456 => x"08",		-- 00d8a0: 084C             MOV.W   R12,R8
						   55457 => x"2C",
						   55458 => x"2C",		-- 00d8a2: 2C48             MOV.W   @R8,R12
						   55459 => x"28",
						   55460 => x"3D",		-- 00d8a4: 3D40             MOV.W   #0x003a,R13
						   55461 => x"20",
						   55462 => x"3A",		-- 00d8a6: 3A00            
						   55463 => x"00",
						   55464 => x"B0",		-- 00d8a8: B012             CALL    #strchr
						   55465 => x"F2",
						   55466 => x"A0",		-- 00d8aa: A0E0            
						   55467 => x"E0",
						   55468 => x"09",		-- 00d8ac: 094C             MOV.W   R12,R9
						   55469 => x"2C",
						   55470 => x"09",		-- 00d8ae: 0993             TST.W   R9
						   55471 => x"73",
						   55472 => x"18",		-- 00d8b0: 1824             JEQ     ($C$L5)
						   55473 => x"04",
						   55474 => x"0A",		-- 00d8b2: 0A49             MOV.W   R9,R10
						   55475 => x"29",
						   55476 => x"2A",		-- 00d8b4: 2A88             SUB.W   @R8,R10
						   55477 => x"68",
						   55478 => x"3A",		-- 00d8b6: 3A90             CMP.W   #0x0009,R10
						   55479 => x"70",
						   55480 => x"09",		-- 00d8b8: 0900            
						   55481 => x"00",
						   55482 => x"01",		-- 00d8ba: 0138             JL      ($C$L4)
						   55483 => x"18",
						   55484 => x"3A",		-- 00d8bc: 3A42             MOV.W   #8,R10
						   55485 => x"22",
						   55486 => x"2D",		-- 00d8be: 2D48             MOV.W   @R8,R13
						   55487 => x"28",
						   55488 => x"0E",		-- 00d8c0: 0E4A             MOV.W   R10,R14
						   55489 => x"2A",
						   55490 => x"0C",		-- 00d8c2: 0C41             MOV.W   SP,R12
						   55491 => x"21",
						   55492 => x"B0",		-- 00d8c4: B012             CALL    #strncpy
						   55493 => x"F2",
						   55494 => x"C8",		-- 00d8c6: C8DE            
						   55495 => x"DE",
						   55496 => x"0F",		-- 00d8c8: 0F41             MOV.W   SP,R15
						   55497 => x"21",
						   55498 => x"0F",		-- 00d8ca: 0F5A             ADD.W   R10,R15
						   55499 => x"3A",
						   55500 => x"CF",		-- 00d8cc: CF43             CLR.B   0x0000(R15)
						   55501 => x"23",
						   55502 => x"00",		-- 00d8ce: 0000            
						   55503 => x"00",
						   55504 => x"0C",		-- 00d8d0: 0C41             MOV.W   SP,R12
						   55505 => x"21",
						   55506 => x"B0",		-- 00d8d2: B012             CALL    #finddevice
						   55507 => x"F2",
						   55508 => x"86",		-- 00d8d4: 86DD            
						   55509 => x"DD",
						   55510 => x"0C",		-- 00d8d6: 0C93             TST.W   R12
						   55511 => x"73",
						   55512 => x"04",		-- 00d8d8: 0424             JEQ     ($C$L5)
						   55513 => x"04",
						   55514 => x"19",		-- 00d8da: 1953             INC.W   R9
						   55515 => x"33",
						   55516 => x"88",		-- 00d8dc: 8849             MOV.W   R9,0x0000(R8)
						   55517 => x"29",
						   55518 => x"00",		-- 00d8de: 0000            
						   55519 => x"00",
						   55520 => x"02",		-- 00d8e0: 023C             JMP     ($C$L6)
						   55521 => x"1C",
						   55522 => x"3C",		-- 00d8e2: 3C40             MOV.W   #0x2078,R12
						   55523 => x"20",
						   55524 => x"78",		-- 00d8e4: 7820            
						   55525 => x"20",
						   55526 => x"31",		-- 00d8e6: 3150             ADD.W   #0x000a,SP
						   55527 => x"30",
						   55528 => x"0A",		-- 00d8e8: 0A00            
						   55529 => x"00",
						   55530 => x"30",		-- 00d8ea: 3040             BR      #__mspabi_func_epilog_3
						   55531 => x"20",
						   55532 => x"9C",		-- 00d8ec: 9CE1            
						   55533 => x"E1",
						   -- Begin: __mspabi_divul
						   -- Begin: __mspabi_remul
						   55534 => x"0A",		-- 00d8ee: 0A12             PUSH    R10
						   55535 => x"F2",
						   55536 => x"09",		-- 00d8f0: 0912             PUSH    R9
						   55537 => x"F2",
						   55538 => x"09",		-- 00d8f2: 0943             CLR.W   R9
						   55539 => x"23",
						   55540 => x"0A",		-- 00d8f4: 0A43             CLR.W   R10
						   55541 => x"23",
						   55542 => x"1B",		-- 00d8f6: 1B43             MOV.W   #1,R11
						   55543 => x"23",
						   55544 => x"0F",		-- 00d8f8: 0F93             TST.W   R15
						   55545 => x"73",
						   55546 => x"04",		-- 00d8fa: 0424             JEQ     (div_loop_lo)
						   55547 => x"04",
						   55548 => x"09",		-- 00d8fc: 094D             MOV.W   R13,R9
						   55549 => x"2D",
						   55550 => x"0D",		-- 00d8fe: 0D4C             MOV.W   R12,R13
						   55551 => x"2C",
						   55552 => x"0C",		-- 00d900: 0C43             CLR.W   R12
						   55553 => x"23",
						   55554 => x"0D",		-- 00d902: 0D3C             JMP     (div_loop_hi)
						   55555 => x"1C",
						   -- Begin: div_loop_lo
						   55556 => x"0C",		-- 00d904: 0C5C             RLA.W   R12
						   55557 => x"3C",
						   55558 => x"0D",		-- 00d906: 0D6D             RLC.W   R13
						   55559 => x"4D",
						   55560 => x"09",		-- 00d908: 0969             RLC.W   R9
						   55561 => x"49",
						   55562 => x"09",		-- 00d90a: 098E             SUB.W   R14,R9
						   55563 => x"6E",
						   55564 => x"04",		-- 00d90c: 0428             JLO     (undo_sub)
						   55565 => x"08",
						   55566 => x"1C",		-- 00d90e: 1CD3             BIS.W   #1,R12
						   55567 => x"B3",
						   55568 => x"0B",		-- 00d910: 0B5B             RLA.W   R11
						   55569 => x"3B",
						   55570 => x"F8",		-- 00d912: F82B             JLO     (div_loop_lo)
						   55571 => x"0B",
						   55572 => x"03",		-- 00d914: 033C             JMP     (process_hi)
						   55573 => x"1C",
						   -- Begin: undo_sub
						   55574 => x"09",		-- 00d916: 095E             ADD.W   R14,R9
						   55575 => x"3E",
						   55576 => x"0B",		-- 00d918: 0B5B             RLA.W   R11
						   55577 => x"3B",
						   55578 => x"F4",		-- 00d91a: F42B             JLO     (div_loop_lo)
						   55579 => x"0B",
						   -- Begin: process_hi
						   55580 => x"1B",		-- 00d91c: 1B43             MOV.W   #1,R11
						   55581 => x"23",
						   -- Begin: div_loop_hi
						   55582 => x"0C",		-- 00d91e: 0C5C             RLA.W   R12
						   55583 => x"3C",
						   55584 => x"0D",		-- 00d920: 0D6D             RLC.W   R13
						   55585 => x"4D",
						   55586 => x"09",		-- 00d922: 0969             RLC.W   R9
						   55587 => x"49",
						   55588 => x"0A",		-- 00d924: 0A6A             RLC.W   R10
						   55589 => x"4A",
						   55590 => x"09",		-- 00d926: 098E             SUB.W   R14,R9
						   55591 => x"6E",
						   55592 => x"0A",		-- 00d928: 0A7F             SUBC.W  R15,R10
						   55593 => x"5F",
						   55594 => x"04",		-- 00d92a: 0428             JLO     (undo_sub_hi)
						   55595 => x"08",
						   55596 => x"1C",		-- 00d92c: 1CD3             BIS.W   #1,R12
						   55597 => x"B3",
						   55598 => x"0B",		-- 00d92e: 0B5B             RLA.W   R11
						   55599 => x"3B",
						   55600 => x"F6",		-- 00d930: F62B             JLO     (div_loop_hi)
						   55601 => x"0B",
						   55602 => x"04",		-- 00d932: 043C             JMP     (div_end)
						   55603 => x"1C",
						   -- Begin: undo_sub_hi
						   55604 => x"09",		-- 00d934: 095E             ADD.W   R14,R9
						   55605 => x"3E",
						   55606 => x"0A",		-- 00d936: 0A6F             ADDC.W  R15,R10
						   55607 => x"4F",
						   55608 => x"0B",		-- 00d938: 0B5B             RLA.W   R11
						   55609 => x"3B",
						   55610 => x"F1",		-- 00d93a: F12B             JLO     (div_loop_hi)
						   55611 => x"0B",
						   -- Begin: div_end
						   55612 => x"0E",		-- 00d93c: 0E49             MOV.W   R9,R14
						   55613 => x"29",
						   55614 => x"0F",		-- 00d93e: 0F4A             MOV.W   R10,R15
						   55615 => x"2A",
						   55616 => x"39",		-- 00d940: 3941             POP.W   R9
						   55617 => x"21",
						   55618 => x"3A",		-- 00d942: 3A41             POP.W   R10
						   55619 => x"21",
						   55620 => x"30",		-- 00d944: 3041             RET     
						   55621 => x"21",
						   -- Begin: atoi
						   55622 => x"0A",		-- 00d946: 0A12             PUSH    R10
						   55623 => x"F2",
						   55624 => x"0B",		-- 00d948: 0B4C             MOV.W   R12,R11
						   55625 => x"2C",
						   55626 => x"0C",		-- 00d94a: 0C43             CLR.W   R12
						   55627 => x"23",
						   55628 => x"0B",		-- 00d94c: 0B3C             JMP     ($C$L3)
						   55629 => x"1C",
						   55630 => x"3D",		-- 00d94e: 3D40             MOV.W   #0x000a,R13
						   55631 => x"20",
						   55632 => x"0A",		-- 00d950: 0A00            
						   55633 => x"00",
						   55634 => x"B0",		-- 00d952: B012             CALL    #__mspabi_mpyi
						   55635 => x"F2",
						   55636 => x"24",		-- 00d954: 24E1            
						   55637 => x"E1",
						   55638 => x"0C",		-- 00d956: 0C5F             ADD.W   R15,R12
						   55639 => x"3F",
						   55640 => x"3C",		-- 00d958: 3C80             SUB.W   #0x0030,R12
						   55641 => x"60",
						   55642 => x"30",		-- 00d95a: 3000            
						   55643 => x"00",
						   55644 => x"1B",		-- 00d95c: 1B53             INC.W   R11
						   55645 => x"33",
						   55646 => x"6F",		-- 00d95e: 6F4B             MOV.B   @R11,R15
						   55647 => x"2B",
						   55648 => x"12",		-- 00d960: 123C             JMP     ($C$L6)
						   55649 => x"1C",
						   55650 => x"1B",		-- 00d962: 1B53             INC.W   R11
						   55651 => x"33",
						   55652 => x"6F",		-- 00d964: 6F4B             MOV.B   @R11,R15
						   55653 => x"2B",
						   55654 => x"4E",		-- 00d966: 4E4F             MOV.B   R15,R14
						   55655 => x"2F",
						   55656 => x"FE",		-- 00d968: FEB2             BIT.B   #8,0x992f(R14)
						   55657 => x"92",
						   55658 => x"2F",		-- 00d96a: 2F99            
						   55659 => x"99",
						   55660 => x"FA",		-- 00d96c: FA23             JNE     ($C$L2)
						   55661 => x"03",
						   55662 => x"4F",		-- 00d96e: 4F4F             MOV.B   R15,R15
						   55663 => x"2F",
						   55664 => x"3F",		-- 00d970: 3F90             CMP.W   #0x002d,R15
						   55665 => x"70",
						   55666 => x"2D",		-- 00d972: 2D00            
						   55667 => x"00",
						   55668 => x"05",		-- 00d974: 0524             JEQ     ($C$L4)
						   55669 => x"04",
						   55670 => x"0A",		-- 00d976: 0A43             CLR.W   R10
						   55671 => x"23",
						   55672 => x"3F",		-- 00d978: 3F90             CMP.W   #0x002b,R15
						   55673 => x"70",
						   55674 => x"2B",		-- 00d97a: 2B00            
						   55675 => x"00",
						   55676 => x"04",		-- 00d97c: 0420             JNE     ($C$L6)
						   55677 => x"00",
						   55678 => x"01",		-- 00d97e: 013C             JMP     ($C$L5)
						   55679 => x"1C",
						   55680 => x"1A",		-- 00d980: 1A43             MOV.W   #1,R10
						   55681 => x"23",
						   55682 => x"1B",		-- 00d982: 1B53             INC.W   R11
						   55683 => x"33",
						   55684 => x"6F",		-- 00d984: 6F4B             MOV.B   @R11,R15
						   55685 => x"2B",
						   55686 => x"EF",		-- 00d986: EFB2             BIT.B   #4,0x992f(R15)
						   55687 => x"92",
						   55688 => x"2F",		-- 00d988: 2F99            
						   55689 => x"99",
						   55690 => x"E1",		-- 00d98a: E123             JNE     ($C$L1)
						   55691 => x"03",
						   55692 => x"0A",		-- 00d98c: 0A93             TST.W   R10
						   55693 => x"73",
						   55694 => x"02",		-- 00d98e: 0224             JEQ     ($C$L7)
						   55695 => x"04",
						   55696 => x"3C",		-- 00d990: 3CE3             INV.W   R12
						   55697 => x"C3",
						   55698 => x"1C",		-- 00d992: 1C53             INC.W   R12
						   55699 => x"33",
						   55700 => x"3A",		-- 00d994: 3A41             POP.W   R10
						   55701 => x"21",
						   55702 => x"30",		-- 00d996: 3041             RET     
						   55703 => x"21",
						   -- Begin: _fcpy
						   55704 => x"0A",		-- 00d998: 0A12             PUSH    R10
						   55705 => x"F2",
						   55706 => x"09",		-- 00d99a: 0912             PUSH    R9
						   55707 => x"F2",
						   55708 => x"08",		-- 00d99c: 0812             PUSH    R8
						   55709 => x"F2",
						   55710 => x"07",		-- 00d99e: 0712             PUSH    R7
						   55711 => x"F2",
						   55712 => x"08",		-- 00d9a0: 084F             MOV.W   R15,R8
						   55713 => x"2F",
						   55714 => x"09",		-- 00d9a2: 094E             MOV.W   R14,R9
						   55715 => x"2E",
						   55716 => x"07",		-- 00d9a4: 074C             MOV.W   R12,R7
						   55717 => x"2C",
						   55718 => x"0D",		-- 00d9a6: 0D59             ADD.W   R9,R13
						   55719 => x"39",
						   55720 => x"1D",		-- 00d9a8: 1D83             DEC.W   R13
						   55721 => x"63",
						   55722 => x"0A",		-- 00d9aa: 0A4D             MOV.W   R13,R10
						   55723 => x"2D",
						   55724 => x"B0",		-- 00d9ac: B012             CALL    #strlen
						   55725 => x"F2",
						   55726 => x"B4",		-- 00d9ae: B4E1            
						   55727 => x"E1",
						   55728 => x"19",		-- 00d9b0: 1983             DEC.W   R9
						   55729 => x"63",
						   55730 => x"09",		-- 00d9b2: 0993             TST.W   R9
						   55731 => x"73",
						   55732 => x"16",		-- 00d9b4: 1638             JL      ($C$L149)
						   55733 => x"18",
						   55734 => x"1E",		-- 00d9b6: 1E43             MOV.W   #1,R14
						   55735 => x"23",
						   55736 => x"0E",		-- 00d9b8: 0E59             ADD.W   R9,R14
						   55737 => x"39",
						   55738 => x"0A",		-- 00d9ba: 0A93             TST.W   R10
						   55739 => x"73",
						   55740 => x"06",		-- 00d9bc: 0638             JL      ($C$L147)
						   55741 => x"18",
						   55742 => x"0A",		-- 00d9be: 0A9C             CMP.W   R12,R10
						   55743 => x"7C",
						   55744 => x"04",		-- 00d9c0: 0434             JGE     ($C$L147)
						   55745 => x"14",
						   55746 => x"0F",		-- 00d9c2: 0F4A             MOV.W   R10,R15
						   55747 => x"2A",
						   55748 => x"0F",		-- 00d9c4: 0F57             ADD.W   R7,R15
						   55749 => x"37",
						   55750 => x"6D",		-- 00d9c6: 6D4F             MOV.B   @R15,R13
						   55751 => x"2F",
						   55752 => x"02",		-- 00d9c8: 023C             JMP     ($C$L148)
						   55753 => x"1C",
						   55754 => x"3D",		-- 00d9ca: 3D40             MOV.W   #0x0030,R13
						   55755 => x"20",
						   55756 => x"30",		-- 00d9cc: 3000            
						   55757 => x"00",
						   55758 => x"2B",		-- 00d9ce: 2B48             MOV.W   @R8,R11
						   55759 => x"28",
						   55760 => x"0F",		-- 00d9d0: 0F4B             MOV.W   R11,R15
						   55761 => x"2B",
						   55762 => x"1F",		-- 00d9d2: 1F83             DEC.W   R15
						   55763 => x"63",
						   55764 => x"88",		-- 00d9d4: 884F             MOV.W   R15,0x0000(R8)
						   55765 => x"2F",
						   55766 => x"00",		-- 00d9d6: 0000            
						   55767 => x"00",
						   55768 => x"CB",		-- 00d9d8: CB4D             MOV.B   R13,0x0000(R11)
						   55769 => x"2D",
						   55770 => x"00",		-- 00d9da: 0000            
						   55771 => x"00",
						   55772 => x"1A",		-- 00d9dc: 1A83             DEC.W   R10
						   55773 => x"63",
						   55774 => x"1E",		-- 00d9de: 1E83             DEC.W   R14
						   55775 => x"63",
						   55776 => x"EC",		-- 00d9e0: EC23             JNE     ($C$L146)
						   55777 => x"03",
						   55778 => x"30",		-- 00d9e2: 3040             BR      #__mspabi_func_epilog_4
						   55779 => x"20",
						   55780 => x"9A",		-- 00d9e4: 9AE1            
						   55781 => x"E1",
						   -- Begin: __mspabi_srli
						   55782 => x"3D",		-- 00d9e6: 3DF0             AND.W   #0x000f,R13
						   55783 => x"D0",
						   55784 => x"0F",		-- 00d9e8: 0F00            
						   55785 => x"00",
						   55786 => x"3D",		-- 00d9ea: 3DE0             XOR.W   #0x000f,R13
						   55787 => x"C0",
						   55788 => x"0F",		-- 00d9ec: 0F00            
						   55789 => x"00",
						   55790 => x"0D",		-- 00d9ee: 0D5D             RLA.W   R13
						   55791 => x"3D",
						   55792 => x"0D",		-- 00d9f0: 0D5D             RLA.W   R13
						   55793 => x"3D",
						   55794 => x"00",		-- 00d9f2: 005D             ADD.W   R13,PC
						   55795 => x"3D",
						   -- Begin: __mspabi_srli_15
						   55796 => x"12",		-- 00d9f4: 12C3             CLRC    
						   55797 => x"A3",
						   55798 => x"0C",		-- 00d9f6: 0C10             RRC     R12
						   55799 => x"F0",
						   -- Begin: __mspabi_srli_14
						   55800 => x"12",		-- 00d9f8: 12C3             CLRC    
						   55801 => x"A3",
						   55802 => x"0C",		-- 00d9fa: 0C10             RRC     R12
						   55803 => x"F0",
						   -- Begin: __mspabi_srli_13
						   55804 => x"12",		-- 00d9fc: 12C3             CLRC    
						   55805 => x"A3",
						   55806 => x"0C",		-- 00d9fe: 0C10             RRC     R12
						   55807 => x"F0",
						   -- Begin: __mspabi_srli_12
						   55808 => x"12",		-- 00da00: 12C3             CLRC    
						   55809 => x"A3",
						   55810 => x"0C",		-- 00da02: 0C10             RRC     R12
						   55811 => x"F0",
						   -- Begin: __mspabi_srli_11
						   55812 => x"12",		-- 00da04: 12C3             CLRC    
						   55813 => x"A3",
						   55814 => x"0C",		-- 00da06: 0C10             RRC     R12
						   55815 => x"F0",
						   -- Begin: __mspabi_srli_10
						   55816 => x"12",		-- 00da08: 12C3             CLRC    
						   55817 => x"A3",
						   55818 => x"0C",		-- 00da0a: 0C10             RRC     R12
						   55819 => x"F0",
						   -- Begin: __mspabi_srli_9
						   55820 => x"12",		-- 00da0c: 12C3             CLRC    
						   55821 => x"A3",
						   55822 => x"0C",		-- 00da0e: 0C10             RRC     R12
						   55823 => x"F0",
						   -- Begin: __mspabi_srli_8
						   55824 => x"12",		-- 00da10: 12C3             CLRC    
						   55825 => x"A3",
						   55826 => x"0C",		-- 00da12: 0C10             RRC     R12
						   55827 => x"F0",
						   -- Begin: __mspabi_srli_7
						   55828 => x"12",		-- 00da14: 12C3             CLRC    
						   55829 => x"A3",
						   55830 => x"0C",		-- 00da16: 0C10             RRC     R12
						   55831 => x"F0",
						   -- Begin: __mspabi_srli_6
						   55832 => x"12",		-- 00da18: 12C3             CLRC    
						   55833 => x"A3",
						   55834 => x"0C",		-- 00da1a: 0C10             RRC     R12
						   55835 => x"F0",
						   -- Begin: __mspabi_srli_5
						   55836 => x"12",		-- 00da1c: 12C3             CLRC    
						   55837 => x"A3",
						   55838 => x"0C",		-- 00da1e: 0C10             RRC     R12
						   55839 => x"F0",
						   -- Begin: __mspabi_srli_4
						   55840 => x"12",		-- 00da20: 12C3             CLRC    
						   55841 => x"A3",
						   55842 => x"0C",		-- 00da22: 0C10             RRC     R12
						   55843 => x"F0",
						   -- Begin: __mspabi_srli_3
						   55844 => x"12",		-- 00da24: 12C3             CLRC    
						   55845 => x"A3",
						   55846 => x"0C",		-- 00da26: 0C10             RRC     R12
						   55847 => x"F0",
						   -- Begin: __mspabi_srli_2
						   55848 => x"12",		-- 00da28: 12C3             CLRC    
						   55849 => x"A3",
						   55850 => x"0C",		-- 00da2a: 0C10             RRC     R12
						   55851 => x"F0",
						   -- Begin: __mspabi_srli_1
						   55852 => x"12",		-- 00da2c: 12C3             CLRC    
						   55853 => x"A3",
						   55854 => x"0C",		-- 00da2e: 0C10             RRC     R12
						   55855 => x"F0",
						   55856 => x"30",		-- 00da30: 3041             RET     
						   55857 => x"21",
						   -- Begin: __mspabi_srall
						   55858 => x"07",		-- 00da32: 0712             PUSH    R7
						   55859 => x"F2",
						   55860 => x"07",		-- 00da34: 074C             MOV.W   R12,R7
						   55861 => x"2C",
						   55862 => x"0D",		-- 00da36: 0D49             MOV.W   R9,R13
						   55863 => x"29",
						   55864 => x"0E",		-- 00da38: 0E4A             MOV.W   R10,R14
						   55865 => x"2A",
						   55866 => x"0F",		-- 00da3a: 0F4B             MOV.W   R11,R15
						   55867 => x"2B",
						   55868 => x"37",		-- 00da3c: 3790             CMP.W   #0x0011,R7
						   55869 => x"70",
						   55870 => x"11",		-- 00da3e: 1100            
						   55871 => x"00",
						   55872 => x"11",		-- 00da40: 1138             JL      ($C$L2)
						   55873 => x"18",
						   55874 => x"0B",		-- 00da42: 0B47             MOV.W   R7,R11
						   55875 => x"27",
						   55876 => x"1B",		-- 00da44: 1B83             DEC.W   R11
						   55877 => x"63",
						   55878 => x"0C",		-- 00da46: 0C4B             MOV.W   R11,R12
						   55879 => x"2B",
						   55880 => x"B0",		-- 00da48: B012             CALL    #__mspabi_srai_4
						   55881 => x"F2",
						   55882 => x"92",		-- 00da4a: 92DE            
						   55883 => x"DE",
						   55884 => x"3B",		-- 00da4c: 3BF0             AND.W   #0xfff0,R11
						   55885 => x"D0",
						   55886 => x"F0",		-- 00da4e: F0FF            
						   55887 => x"FF",
						   55888 => x"07",		-- 00da50: 078B             SUB.W   R11,R7
						   55889 => x"6B",
						   55890 => x"08",		-- 00da52: 084D             MOV.W   R13,R8
						   55891 => x"2D",
						   55892 => x"0D",		-- 00da54: 0D4E             MOV.W   R14,R13
						   55893 => x"2E",
						   55894 => x"0E",		-- 00da56: 0E4F             MOV.W   R15,R14
						   55895 => x"2F",
						   55896 => x"3F",		-- 00da58: 3FB0             BIT.W   #0x8000,R15
						   55897 => x"90",
						   55898 => x"00",		-- 00da5a: 0080            
						   55899 => x"80",
						   55900 => x"0F",		-- 00da5c: 0F7F             SUBC.W  R15,R15
						   55901 => x"5F",
						   55902 => x"3F",		-- 00da5e: 3FE3             INV.W   R15
						   55903 => x"C3",
						   55904 => x"1C",		-- 00da60: 1C83             DEC.W   R12
						   55905 => x"63",
						   55906 => x"F7",		-- 00da62: F723             JNE     ($C$L1)
						   55907 => x"03",
						   55908 => x"17",		-- 00da64: 1793             CMP.W   #1,R7
						   55909 => x"73",
						   55910 => x"07",		-- 00da66: 0738             JL      ($C$L4)
						   55911 => x"18",
						   55912 => x"0C",		-- 00da68: 0C47             MOV.W   R7,R12
						   55913 => x"27",
						   55914 => x"0F",		-- 00da6a: 0F11             RRA     R15
						   55915 => x"F1",
						   55916 => x"0E",		-- 00da6c: 0E10             RRC     R14
						   55917 => x"F0",
						   55918 => x"0D",		-- 00da6e: 0D10             RRC     R13
						   55919 => x"F0",
						   55920 => x"08",		-- 00da70: 0810             RRC     R8
						   55921 => x"F0",
						   55922 => x"1C",		-- 00da72: 1C83             DEC.W   R12
						   55923 => x"63",
						   55924 => x"FA",		-- 00da74: FA23             JNE     ($C$L3)
						   55925 => x"03",
						   55926 => x"0C",		-- 00da76: 0C48             MOV.W   R8,R12
						   55927 => x"28",
						   55928 => x"37",		-- 00da78: 3741             POP.W   R7
						   55929 => x"21",
						   55930 => x"30",		-- 00da7a: 3041             RET     
						   55931 => x"21",
						   -- Begin: close
						   55932 => x"0A",		-- 00da7c: 0A12             PUSH    R10
						   55933 => x"F2",
						   55934 => x"0A",		-- 00da7e: 0A4C             MOV.W   R12,R10
						   55935 => x"2C",
						   55936 => x"0A",		-- 00da80: 0A93             TST.W   R10
						   55937 => x"73",
						   55938 => x"03",		-- 00da82: 0338             JL      ($C$L1)
						   55939 => x"18",
						   55940 => x"3A",		-- 00da84: 3A90             CMP.W   #0x000a,R10
						   55941 => x"70",
						   55942 => x"0A",		-- 00da86: 0A00            
						   55943 => x"00",
						   55944 => x"02",		-- 00da88: 0238             JL      ($C$L2)
						   55945 => x"18",
						   55946 => x"3A",		-- 00da8a: 3A43             MOV.W   #-1,R10
						   55947 => x"23",
						   55948 => x"19",		-- 00da8c: 193C             JMP     ($C$L6)
						   55949 => x"1C",
						   55950 => x"92",		-- 00da8e: 9212             CALL    &_lock
						   55951 => x"F2",
						   55952 => x"F2",		-- 00da90: F220            
						   55953 => x"20",
						   55954 => x"0A",		-- 00da92: 0A5A             RLA.W   R10
						   55955 => x"3A",
						   55956 => x"0A",		-- 00da94: 0A5A             RLA.W   R10
						   55957 => x"3A",
						   55958 => x"3A",		-- 00da96: 3A50             ADD.W   #0x20c6,R10
						   55959 => x"30",
						   55960 => x"C6",		-- 00da98: C620            
						   55961 => x"20",
						   55962 => x"2F",		-- 00da9a: 2F4A             MOV.W   @R10,R15
						   55963 => x"2A",
						   55964 => x"0F",		-- 00da9c: 0F93             TST.W   R15
						   55965 => x"73",
						   55966 => x"02",		-- 00da9e: 0220             JNE     ($C$L3)
						   55967 => x"00",
						   55968 => x"3A",		-- 00daa0: 3A43             MOV.W   #-1,R10
						   55969 => x"23",
						   55970 => x"0C",		-- 00daa2: 0C3C             JMP     ($C$L5)
						   55971 => x"1C",
						   55972 => x"1C",		-- 00daa4: 1C4A             MOV.W   0x0002(R10),R12
						   55973 => x"2A",
						   55974 => x"02",		-- 00daa6: 0200            
						   55975 => x"00",
						   55976 => x"9F",		-- 00daa8: 9F12             CALL    0x000e(R15)
						   55977 => x"F2",
						   55978 => x"0E",		-- 00daaa: 0E00            
						   55979 => x"00",
						   55980 => x"3C",		-- 00daac: 3C93             CMP.W   #-1,R12
						   55981 => x"73",
						   55982 => x"05",		-- 00daae: 0524             JEQ     ($C$L4)
						   55983 => x"04",
						   55984 => x"2F",		-- 00dab0: 2F4A             MOV.W   @R10,R15
						   55985 => x"2A",
						   55986 => x"9F",		-- 00dab2: 9FC3             BIC.W   #1,0x000a(R15)
						   55987 => x"A3",
						   55988 => x"0A",		-- 00dab4: 0A00            
						   55989 => x"00",
						   55990 => x"8A",		-- 00dab6: 8A43             CLR.W   0x0000(R10)
						   55991 => x"23",
						   55992 => x"00",		-- 00dab8: 0000            
						   55993 => x"00",
						   55994 => x"0A",		-- 00daba: 0A4C             MOV.W   R12,R10
						   55995 => x"2C",
						   55996 => x"92",		-- 00dabc: 9212             CALL    &_unlock
						   55997 => x"F2",
						   55998 => x"F4",		-- 00dabe: F420            
						   55999 => x"20",
						   56000 => x"0C",		-- 00dac0: 0C4A             MOV.W   R10,R12
						   56001 => x"2A",
						   56002 => x"3A",		-- 00dac2: 3A41             POP.W   R10
						   56003 => x"21",
						   56004 => x"30",		-- 00dac4: 3041             RET     
						   56005 => x"21",
						   -- Begin: __mspabi_srlll
						   56006 => x"07",		-- 00dac6: 0712             PUSH    R7
						   56007 => x"F2",
						   56008 => x"07",		-- 00dac8: 074C             MOV.W   R12,R7
						   56009 => x"2C",
						   56010 => x"0D",		-- 00daca: 0D49             MOV.W   R9,R13
						   56011 => x"29",
						   56012 => x"0E",		-- 00dacc: 0E4A             MOV.W   R10,R14
						   56013 => x"2A",
						   56014 => x"0F",		-- 00dace: 0F4B             MOV.W   R11,R15
						   56015 => x"2B",
						   56016 => x"37",		-- 00dad0: 3790             CMP.W   #0x0011,R7
						   56017 => x"70",
						   56018 => x"11",		-- 00dad2: 1100            
						   56019 => x"00",
						   56020 => x"0E",		-- 00dad4: 0E38             JL      ($C$L2)
						   56021 => x"18",
						   56022 => x"0B",		-- 00dad6: 0B47             MOV.W   R7,R11
						   56023 => x"27",
						   56024 => x"1B",		-- 00dad8: 1B83             DEC.W   R11
						   56025 => x"63",
						   56026 => x"0C",		-- 00dada: 0C4B             MOV.W   R11,R12
						   56027 => x"2B",
						   56028 => x"B0",		-- 00dadc: B012             CALL    #__mspabi_srai_4
						   56029 => x"F2",
						   56030 => x"92",		-- 00dade: 92DE            
						   56031 => x"DE",
						   56032 => x"3B",		-- 00dae0: 3BF0             AND.W   #0xfff0,R11
						   56033 => x"D0",
						   56034 => x"F0",		-- 00dae2: F0FF            
						   56035 => x"FF",
						   56036 => x"07",		-- 00dae4: 078B             SUB.W   R11,R7
						   56037 => x"6B",
						   56038 => x"08",		-- 00dae6: 084D             MOV.W   R13,R8
						   56039 => x"2D",
						   56040 => x"0D",		-- 00dae8: 0D4E             MOV.W   R14,R13
						   56041 => x"2E",
						   56042 => x"0E",		-- 00daea: 0E4F             MOV.W   R15,R14
						   56043 => x"2F",
						   56044 => x"0F",		-- 00daec: 0F43             CLR.W   R15
						   56045 => x"23",
						   56046 => x"1C",		-- 00daee: 1C83             DEC.W   R12
						   56047 => x"63",
						   56048 => x"FA",		-- 00daf0: FA23             JNE     ($C$L1)
						   56049 => x"03",
						   56050 => x"17",		-- 00daf2: 1793             CMP.W   #1,R7
						   56051 => x"73",
						   56052 => x"08",		-- 00daf4: 0838             JL      ($C$L4)
						   56053 => x"18",
						   56054 => x"0C",		-- 00daf6: 0C47             MOV.W   R7,R12
						   56055 => x"27",
						   56056 => x"12",		-- 00daf8: 12C3             CLRC    
						   56057 => x"A3",
						   56058 => x"0F",		-- 00dafa: 0F10             RRC     R15
						   56059 => x"F0",
						   56060 => x"0E",		-- 00dafc: 0E10             RRC     R14
						   56061 => x"F0",
						   56062 => x"0D",		-- 00dafe: 0D10             RRC     R13
						   56063 => x"F0",
						   56064 => x"08",		-- 00db00: 0810             RRC     R8
						   56065 => x"F0",
						   56066 => x"1C",		-- 00db02: 1C83             DEC.W   R12
						   56067 => x"63",
						   56068 => x"F9",		-- 00db04: F923             JNE     ($C$L3)
						   56069 => x"03",
						   56070 => x"0C",		-- 00db06: 0C48             MOV.W   R8,R12
						   56071 => x"28",
						   56072 => x"37",		-- 00db08: 3741             POP.W   R7
						   56073 => x"21",
						   56074 => x"30",		-- 00db0a: 3041             RET     
						   56075 => x"21",
						   -- Begin: HOSTclose
						   56076 => x"0A",		-- 00db0c: 0A12             PUSH    R10
						   56077 => x"F2",
						   56078 => x"0A",		-- 00db0e: 0A4C             MOV.W   R12,R10
						   56079 => x"2C",
						   56080 => x"92",		-- 00db10: 9212             CALL    &_lock
						   56081 => x"F2",
						   56082 => x"F2",		-- 00db12: F220            
						   56083 => x"20",
						   56084 => x"C2",		-- 00db14: C24A             MOV.B   R10,&parmbuf
						   56085 => x"2A",
						   56086 => x"9E",		-- 00db16: 9E21            
						   56087 => x"21",
						   56088 => x"8A",		-- 00db18: 8A10             SWPB    R10
						   56089 => x"F0",
						   56090 => x"8A",		-- 00db1a: 8A11             SXT     R10
						   56091 => x"F1",
						   56092 => x"C2",		-- 00db1c: C24A             MOV.B   R10,&0x219f
						   56093 => x"2A",
						   56094 => x"9F",		-- 00db1e: 9F21            
						   56095 => x"21",
						   56096 => x"7C",		-- 00db20: 7C40             MOV.B   #0x00f1,R12
						   56097 => x"20",
						   56098 => x"F1",		-- 00db22: F100            
						   56099 => x"00",
						   56100 => x"3D",		-- 00db24: 3D40             MOV.W   #0x219e,R13
						   56101 => x"20",
						   56102 => x"9E",		-- 00db26: 9E21            
						   56103 => x"21",
						   56104 => x"0E",		-- 00db28: 0E43             CLR.W   R14
						   56105 => x"23",
						   56106 => x"0F",		-- 00db2a: 0F43             CLR.W   R15
						   56107 => x"23",
						   56108 => x"B0",		-- 00db2c: B012             CALL    #__TI_writemsg
						   56109 => x"F2",
						   56110 => x"BA",		-- 00db2e: BADD            
						   56111 => x"DD",
						   56112 => x"3C",		-- 00db30: 3C40             MOV.W   #0x219e,R12
						   56113 => x"20",
						   56114 => x"9E",		-- 00db32: 9E21            
						   56115 => x"21",
						   56116 => x"0D",		-- 00db34: 0D43             CLR.W   R13
						   56117 => x"23",
						   56118 => x"B0",		-- 00db36: B012             CALL    #__TI_readmsg
						   56119 => x"F2",
						   56120 => x"44",		-- 00db38: 44DE            
						   56121 => x"DE",
						   56122 => x"5F",		-- 00db3a: 5F42             MOV.B   &parmbuf,R15
						   56123 => x"22",
						   56124 => x"9E",		-- 00db3c: 9E21            
						   56125 => x"21",
						   56126 => x"5A",		-- 00db3e: 5A42             MOV.B   &0x219f,R10
						   56127 => x"22",
						   56128 => x"9F",		-- 00db40: 9F21            
						   56129 => x"21",
						   56130 => x"8A",		-- 00db42: 8A10             SWPB    R10
						   56131 => x"F0",
						   56132 => x"0A",		-- 00db44: 0A5F             ADD.W   R15,R10
						   56133 => x"3F",
						   56134 => x"92",		-- 00db46: 9212             CALL    &_unlock
						   56135 => x"F2",
						   56136 => x"F4",		-- 00db48: F420            
						   56137 => x"20",
						   56138 => x"0C",		-- 00db4a: 0C4A             MOV.W   R10,R12
						   56139 => x"2A",
						   56140 => x"3A",		-- 00db4c: 3A41             POP.W   R10
						   56141 => x"21",
						   56142 => x"30",		-- 00db4e: 3041             RET     
						   56143 => x"21",
						   -- Begin: __mspabi_sllll
						   56144 => x"07",		-- 00db50: 0712             PUSH    R7
						   56145 => x"F2",
						   56146 => x"07",		-- 00db52: 074C             MOV.W   R12,R7
						   56147 => x"2C",
						   56148 => x"0D",		-- 00db54: 0D49             MOV.W   R9,R13
						   56149 => x"29",
						   56150 => x"0E",		-- 00db56: 0E4A             MOV.W   R10,R14
						   56151 => x"2A",
						   56152 => x"0F",		-- 00db58: 0F4B             MOV.W   R11,R15
						   56153 => x"2B",
						   56154 => x"37",		-- 00db5a: 3790             CMP.W   #0x0011,R7
						   56155 => x"70",
						   56156 => x"11",		-- 00db5c: 1100            
						   56157 => x"00",
						   56158 => x"0E",		-- 00db5e: 0E38             JL      ($C$L2)
						   56159 => x"18",
						   56160 => x"0F",		-- 00db60: 0F47             MOV.W   R7,R15
						   56161 => x"27",
						   56162 => x"1F",		-- 00db62: 1F83             DEC.W   R15
						   56163 => x"63",
						   56164 => x"0C",		-- 00db64: 0C4F             MOV.W   R15,R12
						   56165 => x"2F",
						   56166 => x"B0",		-- 00db66: B012             CALL    #__mspabi_srai_4
						   56167 => x"F2",
						   56168 => x"92",		-- 00db68: 92DE            
						   56169 => x"DE",
						   56170 => x"3F",		-- 00db6a: 3FF0             AND.W   #0xfff0,R15
						   56171 => x"D0",
						   56172 => x"F0",		-- 00db6c: F0FF            
						   56173 => x"FF",
						   56174 => x"07",		-- 00db6e: 078F             SUB.W   R15,R7
						   56175 => x"6F",
						   56176 => x"0F",		-- 00db70: 0F4E             MOV.W   R14,R15
						   56177 => x"2E",
						   56178 => x"0E",		-- 00db72: 0E4D             MOV.W   R13,R14
						   56179 => x"2D",
						   56180 => x"0D",		-- 00db74: 0D48             MOV.W   R8,R13
						   56181 => x"28",
						   56182 => x"08",		-- 00db76: 0843             CLR.W   R8
						   56183 => x"23",
						   56184 => x"1C",		-- 00db78: 1C83             DEC.W   R12
						   56185 => x"63",
						   56186 => x"FA",		-- 00db7a: FA23             JNE     ($C$L1)
						   56187 => x"03",
						   56188 => x"17",		-- 00db7c: 1793             CMP.W   #1,R7
						   56189 => x"73",
						   56190 => x"07",		-- 00db7e: 0738             JL      ($C$L4)
						   56191 => x"18",
						   56192 => x"0C",		-- 00db80: 0C47             MOV.W   R7,R12
						   56193 => x"27",
						   56194 => x"08",		-- 00db82: 0858             RLA.W   R8
						   56195 => x"38",
						   56196 => x"0D",		-- 00db84: 0D6D             RLC.W   R13
						   56197 => x"4D",
						   56198 => x"0E",		-- 00db86: 0E6E             RLC.W   R14
						   56199 => x"4E",
						   56200 => x"0F",		-- 00db88: 0F6F             RLC.W   R15
						   56201 => x"4F",
						   56202 => x"1C",		-- 00db8a: 1C83             DEC.W   R12
						   56203 => x"63",
						   56204 => x"FA",		-- 00db8c: FA23             JNE     ($C$L3)
						   56205 => x"03",
						   56206 => x"0C",		-- 00db8e: 0C48             MOV.W   R8,R12
						   56207 => x"28",
						   56208 => x"37",		-- 00db90: 3741             POP.W   R7
						   56209 => x"21",
						   56210 => x"30",		-- 00db92: 3041             RET     
						   56211 => x"21",
						   -- Begin: exit
						   56212 => x"0A",		-- 00db94: 0A12             PUSH    R10
						   56213 => x"F2",
						   56214 => x"0A",		-- 00db96: 0A4C             MOV.W   R12,R10
						   56215 => x"2C",
						   56216 => x"82",		-- 00db98: 8293             TST.W   &__TI_enable_exit_profile_output
						   56217 => x"73",
						   56218 => x"FA",		-- 00db9a: FA20            
						   56219 => x"20",
						   56220 => x"0A",		-- 00db9c: 0A24             JEQ     ($C$L3)
						   56221 => x"04",
						   56222 => x"3E",		-- 00db9e: 3E40             MOV.W   #0xffff,R14
						   56223 => x"20",
						   56224 => x"FF",		-- 00dba0: FFFF            
						   56225 => x"FF",
						   56226 => x"3F",		-- 00dba2: 3F40             MOV.W   #0xffff,R15
						   56227 => x"20",
						   56228 => x"FF",		-- 00dba4: FFFF            
						   56229 => x"FF",
						   56230 => x"3F",		-- 00dba6: 3F93             CMP.W   #-1,R15
						   56231 => x"73",
						   56232 => x"02",		-- 00dba8: 0220             JNE     ($C$L2)
						   56233 => x"00",
						   56234 => x"3E",		-- 00dbaa: 3E93             CMP.W   #-1,R14
						   56235 => x"73",
						   56236 => x"02",		-- 00dbac: 0224             JEQ     ($C$L3)
						   56237 => x"04",
						   56238 => x"B0",		-- 00dbae: B012             CALL    #0xffff
						   56239 => x"F2",
						   56240 => x"FF",		-- 00dbb0: FFFF            
						   56241 => x"FF",
						   56242 => x"92",		-- 00dbb2: 9212             CALL    &_lock
						   56243 => x"F2",
						   56244 => x"F2",		-- 00dbb4: F220            
						   56245 => x"20",
						   56246 => x"82",		-- 00dbb6: 8293             TST.W   &__TI_dtors_ptr
						   56247 => x"73",
						   56248 => x"F0",		-- 00dbb8: F020            
						   56249 => x"20",
						   56250 => x"03",		-- 00dbba: 0324             JEQ     ($C$L4)
						   56251 => x"04",
						   56252 => x"0C",		-- 00dbbc: 0C4A             MOV.W   R10,R12
						   56253 => x"2A",
						   56254 => x"92",		-- 00dbbe: 9212             CALL    &__TI_dtors_ptr
						   56255 => x"F2",
						   56256 => x"F0",		-- 00dbc0: F020            
						   56257 => x"20",
						   56258 => x"82",		-- 00dbc2: 8293             TST.W   &__TI_cleanup_ptr
						   56259 => x"73",
						   56260 => x"EE",		-- 00dbc4: EE20            
						   56261 => x"20",
						   56262 => x"02",		-- 00dbc6: 0224             JEQ     ($C$L5)
						   56263 => x"04",
						   56264 => x"92",		-- 00dbc8: 9212             CALL    &__TI_cleanup_ptr
						   56265 => x"F2",
						   56266 => x"EE",		-- 00dbca: EE20            
						   56267 => x"20",
						   56268 => x"92",		-- 00dbcc: 9212             CALL    &_unlock
						   56269 => x"F2",
						   56270 => x"F4",		-- 00dbce: F420            
						   56271 => x"20",
						   56272 => x"B0",		-- 00dbd0: B012             CALL    #abort
						   56273 => x"F2",
						   56274 => x"F2",		-- 00dbd2: F2E1            
						   56275 => x"E1",
						   56276 => x"3A",		-- 00dbd4: 3A41             POP.W   R10
						   56277 => x"21",
						   56278 => x"30",		-- 00dbd6: 3041             RET     
						   56279 => x"21",
						   -- Begin: __TI_auto_init_nobinit_nopinit
						   56280 => x"0A",		-- 00dbd8: 0A12             PUSH    R10
						   56281 => x"F2",
						   56282 => x"09",		-- 00dbda: 0912             PUSH    R9
						   56283 => x"F2",
						   56284 => x"3F",		-- 00dbdc: 3F40             MOV.W   #0x8502,R15
						   56285 => x"20",
						   56286 => x"02",		-- 00dbde: 0285            
						   56287 => x"85",
						   56288 => x"3F",		-- 00dbe0: 3F90             CMP.W   #0x8508,R15
						   56289 => x"70",
						   56290 => x"08",		-- 00dbe2: 0885            
						   56291 => x"85",
						   56292 => x"16",		-- 00dbe4: 1624             JEQ     ($C$L22)
						   56293 => x"04",
						   56294 => x"3F",		-- 00dbe6: 3F40             MOV.W   #0x850c,R15
						   56295 => x"20",
						   56296 => x"0C",		-- 00dbe8: 0C85            
						   56297 => x"85",
						   56298 => x"3F",		-- 00dbea: 3F90             CMP.W   #0x8514,R15
						   56299 => x"70",
						   56300 => x"14",		-- 00dbec: 1485            
						   56301 => x"85",
						   56302 => x"11",		-- 00dbee: 1124             JEQ     ($C$L22)
						   56303 => x"04",
						   56304 => x"3A",		-- 00dbf0: 3A40             MOV.W   #0x8514,R10
						   56305 => x"20",
						   56306 => x"14",		-- 00dbf2: 1485            
						   56307 => x"85",
						   56308 => x"3A",		-- 00dbf4: 3A80             SUB.W   #0x850c,R10
						   56309 => x"60",
						   56310 => x"0C",		-- 00dbf6: 0C85            
						   56311 => x"85",
						   56312 => x"0A",		-- 00dbf8: 0A11             RRA     R10
						   56313 => x"F1",
						   56314 => x"0A",		-- 00dbfa: 0A11             RRA     R10
						   56315 => x"F1",
						   56316 => x"39",		-- 00dbfc: 3940             MOV.W   #0x850c,R9
						   56317 => x"20",
						   56318 => x"0C",		-- 00dbfe: 0C85            
						   56319 => x"85",
						   56320 => x"3C",		-- 00dc00: 3C49             MOV.W   @R9+,R12
						   56321 => x"29",
						   56322 => x"7F",		-- 00dc02: 7F4C             MOV.B   @R12+,R15
						   56323 => x"2C",
						   56324 => x"0F",		-- 00dc04: 0F5F             RLA.W   R15
						   56325 => x"3F",
						   56326 => x"1F",		-- 00dc06: 1F4F             MOV.W   0x8502(R15),R15
						   56327 => x"2F",
						   56328 => x"02",		-- 00dc08: 0285            
						   56329 => x"85",
						   56330 => x"3D",		-- 00dc0a: 3D49             MOV.W   @R9+,R13
						   56331 => x"29",
						   56332 => x"8F",		-- 00dc0c: 8F12             CALL    R15
						   56333 => x"F2",
						   56334 => x"1A",		-- 00dc0e: 1A83             DEC.W   R10
						   56335 => x"63",
						   56336 => x"F7",		-- 00dc10: F723             JNE     ($C$L21)
						   56337 => x"03",
						   56338 => x"B0",		-- 00dc12: B012             CALL    #_system_post_cinit
						   56339 => x"F2",
						   56340 => x"02",		-- 00dc14: 02E2            
						   56341 => x"E2",
						   56342 => x"30",		-- 00dc16: 3040             BR      #__mspabi_func_epilog_2
						   56343 => x"20",
						   56344 => x"9E",		-- 00dc18: 9EE1            
						   56345 => x"E1",
						   -- Begin: HOSTunlink
						   56346 => x"0A",		-- 00dc1a: 0A12             PUSH    R10
						   56347 => x"F2",
						   56348 => x"0A",		-- 00dc1c: 0A4C             MOV.W   R12,R10
						   56349 => x"2C",
						   56350 => x"92",		-- 00dc1e: 9212             CALL    &_lock
						   56351 => x"F2",
						   56352 => x"F2",		-- 00dc20: F220            
						   56353 => x"20",
						   56354 => x"0C",		-- 00dc22: 0C4A             MOV.W   R10,R12
						   56355 => x"2A",
						   56356 => x"B0",		-- 00dc24: B012             CALL    #strlen
						   56357 => x"F2",
						   56358 => x"B4",		-- 00dc26: B4E1            
						   56359 => x"E1",
						   56360 => x"1F",		-- 00dc28: 1F43             MOV.W   #1,R15
						   56361 => x"23",
						   56362 => x"0F",		-- 00dc2a: 0F5C             ADD.W   R12,R15
						   56363 => x"3C",
						   56364 => x"7C",		-- 00dc2c: 7C40             MOV.B   #0x00f5,R12
						   56365 => x"20",
						   56366 => x"F5",		-- 00dc2e: F500            
						   56367 => x"00",
						   56368 => x"3D",		-- 00dc30: 3D40             MOV.W   #0x219e,R13
						   56369 => x"20",
						   56370 => x"9E",		-- 00dc32: 9E21            
						   56371 => x"21",
						   56372 => x"0E",		-- 00dc34: 0E4A             MOV.W   R10,R14
						   56373 => x"2A",
						   56374 => x"B0",		-- 00dc36: B012             CALL    #__TI_writemsg
						   56375 => x"F2",
						   56376 => x"BA",		-- 00dc38: BADD            
						   56377 => x"DD",
						   56378 => x"3C",		-- 00dc3a: 3C40             MOV.W   #0x219e,R12
						   56379 => x"20",
						   56380 => x"9E",		-- 00dc3c: 9E21            
						   56381 => x"21",
						   56382 => x"0D",		-- 00dc3e: 0D43             CLR.W   R13
						   56383 => x"23",
						   56384 => x"B0",		-- 00dc40: B012             CALL    #__TI_readmsg
						   56385 => x"F2",
						   56386 => x"44",		-- 00dc42: 44DE            
						   56387 => x"DE",
						   56388 => x"5F",		-- 00dc44: 5F42             MOV.B   &parmbuf,R15
						   56389 => x"22",
						   56390 => x"9E",		-- 00dc46: 9E21            
						   56391 => x"21",
						   56392 => x"5A",		-- 00dc48: 5A42             MOV.B   &0x219f,R10
						   56393 => x"22",
						   56394 => x"9F",		-- 00dc4a: 9F21            
						   56395 => x"21",
						   56396 => x"8A",		-- 00dc4c: 8A10             SWPB    R10
						   56397 => x"F0",
						   56398 => x"0A",		-- 00dc4e: 0A5F             ADD.W   R15,R10
						   56399 => x"3F",
						   56400 => x"92",		-- 00dc50: 9212             CALL    &_unlock
						   56401 => x"F2",
						   56402 => x"F4",		-- 00dc52: F420            
						   56403 => x"20",
						   56404 => x"0C",		-- 00dc54: 0C4A             MOV.W   R10,R12
						   56405 => x"2A",
						   56406 => x"3A",		-- 00dc56: 3A41             POP.W   R10
						   56407 => x"21",
						   56408 => x"30",		-- 00dc58: 3041             RET     
						   56409 => x"21",
						   -- Begin: __mspabi_divli
						   -- Begin: __mspabi_remli
						   56410 => x"0A",		-- 00dc5a: 0A12             PUSH    R10
						   56411 => x"F2",
						   56412 => x"0A",		-- 00dc5c: 0A43             CLR.W   R10
						   56413 => x"23",
						   56414 => x"0F",		-- 00dc5e: 0F93             TST.W   R15
						   56415 => x"73",
						   56416 => x"05",		-- 00dc60: 0534             JGE     (dvd_sign)
						   56417 => x"14",
						   56418 => x"3E",		-- 00dc62: 3EE3             INV.W   R14
						   56419 => x"C3",
						   56420 => x"3F",		-- 00dc64: 3FE3             INV.W   R15
						   56421 => x"C3",
						   56422 => x"1E",		-- 00dc66: 1E53             INC.W   R14
						   56423 => x"33",
						   56424 => x"0F",		-- 00dc68: 0F63             ADC.W   R15
						   56425 => x"43",
						   56426 => x"1A",		-- 00dc6a: 1AD3             BIS.W   #1,R10
						   56427 => x"B3",
						   -- Begin: dvd_sign
						   56428 => x"0D",		-- 00dc6c: 0D93             TST.W   R13
						   56429 => x"73",
						   56430 => x"05",		-- 00dc6e: 0534             JGE     (perform_divide)
						   56431 => x"14",
						   56432 => x"3C",		-- 00dc70: 3CE3             INV.W   R12
						   56433 => x"C3",
						   56434 => x"3D",		-- 00dc72: 3DE3             INV.W   R13
						   56435 => x"C3",
						   56436 => x"1C",		-- 00dc74: 1C53             INC.W   R12
						   56437 => x"33",
						   56438 => x"0D",		-- 00dc76: 0D63             ADC.W   R13
						   56439 => x"43",
						   56440 => x"3A",		-- 00dc78: 3AE3             INV.W   R10
						   56441 => x"C3",
						   -- Begin: perform_divide
						   56442 => x"B0",		-- 00dc7a: B012             CALL    #__mspabi_divul
						   56443 => x"F2",
						   56444 => x"EE",		-- 00dc7c: EED8            
						   56445 => x"D8",
						   56446 => x"1A",		-- 00dc7e: 1AB3             BIT.W   #1,R10
						   56447 => x"93",
						   56448 => x"04",		-- 00dc80: 0424             JEQ     (rem_sign)
						   56449 => x"04",
						   56450 => x"3C",		-- 00dc82: 3CE3             INV.W   R12
						   56451 => x"C3",
						   56452 => x"3D",		-- 00dc84: 3DE3             INV.W   R13
						   56453 => x"C3",
						   56454 => x"1C",		-- 00dc86: 1C53             INC.W   R12
						   56455 => x"33",
						   56456 => x"0D",		-- 00dc88: 0D63             ADC.W   R13
						   56457 => x"43",
						   -- Begin: rem_sign
						   56458 => x"2A",		-- 00dc8a: 2AB3             BIT.W   #2,R10
						   56459 => x"93",
						   56460 => x"04",		-- 00dc8c: 0424             JEQ     (div_exit)
						   56461 => x"04",
						   56462 => x"3E",		-- 00dc8e: 3EE3             INV.W   R14
						   56463 => x"C3",
						   56464 => x"3F",		-- 00dc90: 3FE3             INV.W   R15
						   56465 => x"C3",
						   56466 => x"1E",		-- 00dc92: 1E53             INC.W   R14
						   56467 => x"33",
						   56468 => x"0F",		-- 00dc94: 0F63             ADC.W   R15
						   56469 => x"43",
						   -- Begin: div_exit
						   56470 => x"3A",		-- 00dc96: 3A41             POP.W   R10
						   56471 => x"21",
						   56472 => x"30",		-- 00dc98: 3041             RET     
						   56473 => x"21",
						   -- Begin: __mspabi_sral_15
						   56474 => x"0D",		-- 00dc9a: 0D11             RRA     R13
						   56475 => x"F1",
						   56476 => x"0C",		-- 00dc9c: 0C10             RRC     R12
						   56477 => x"F0",
						   -- Begin: __mspabi_sral_14
						   56478 => x"0D",		-- 00dc9e: 0D11             RRA     R13
						   56479 => x"F1",
						   56480 => x"0C",		-- 00dca0: 0C10             RRC     R12
						   56481 => x"F0",
						   -- Begin: __mspabi_sral_13
						   56482 => x"0D",		-- 00dca2: 0D11             RRA     R13
						   56483 => x"F1",
						   56484 => x"0C",		-- 00dca4: 0C10             RRC     R12
						   56485 => x"F0",
						   -- Begin: __mspabi_sral_12
						   56486 => x"0D",		-- 00dca6: 0D11             RRA     R13
						   56487 => x"F1",
						   56488 => x"0C",		-- 00dca8: 0C10             RRC     R12
						   56489 => x"F0",
						   -- Begin: __mspabi_sral_11
						   56490 => x"0D",		-- 00dcaa: 0D11             RRA     R13
						   56491 => x"F1",
						   56492 => x"0C",		-- 00dcac: 0C10             RRC     R12
						   56493 => x"F0",
						   -- Begin: __mspabi_sral_10
						   56494 => x"0D",		-- 00dcae: 0D11             RRA     R13
						   56495 => x"F1",
						   56496 => x"0C",		-- 00dcb0: 0C10             RRC     R12
						   56497 => x"F0",
						   -- Begin: __mspabi_sral_9
						   56498 => x"0D",		-- 00dcb2: 0D11             RRA     R13
						   56499 => x"F1",
						   56500 => x"0C",		-- 00dcb4: 0C10             RRC     R12
						   56501 => x"F0",
						   -- Begin: __mspabi_sral_8
						   56502 => x"0D",		-- 00dcb6: 0D11             RRA     R13
						   56503 => x"F1",
						   56504 => x"0C",		-- 00dcb8: 0C10             RRC     R12
						   56505 => x"F0",
						   -- Begin: __mspabi_sral_7
						   56506 => x"0D",		-- 00dcba: 0D11             RRA     R13
						   56507 => x"F1",
						   56508 => x"0C",		-- 00dcbc: 0C10             RRC     R12
						   56509 => x"F0",
						   -- Begin: __mspabi_sral_6
						   56510 => x"0D",		-- 00dcbe: 0D11             RRA     R13
						   56511 => x"F1",
						   56512 => x"0C",		-- 00dcc0: 0C10             RRC     R12
						   56513 => x"F0",
						   -- Begin: __mspabi_sral_5
						   56514 => x"0D",		-- 00dcc2: 0D11             RRA     R13
						   56515 => x"F1",
						   56516 => x"0C",		-- 00dcc4: 0C10             RRC     R12
						   56517 => x"F0",
						   -- Begin: __mspabi_sral_4
						   56518 => x"0D",		-- 00dcc6: 0D11             RRA     R13
						   56519 => x"F1",
						   56520 => x"0C",		-- 00dcc8: 0C10             RRC     R12
						   56521 => x"F0",
						   -- Begin: __mspabi_sral_3
						   56522 => x"0D",		-- 00dcca: 0D11             RRA     R13
						   56523 => x"F1",
						   56524 => x"0C",		-- 00dccc: 0C10             RRC     R12
						   56525 => x"F0",
						   -- Begin: __mspabi_sral_2
						   56526 => x"0D",		-- 00dcce: 0D11             RRA     R13
						   56527 => x"F1",
						   56528 => x"0C",		-- 00dcd0: 0C10             RRC     R12
						   56529 => x"F0",
						   -- Begin: __mspabi_sral_1
						   56530 => x"0D",		-- 00dcd2: 0D11             RRA     R13
						   56531 => x"F1",
						   56532 => x"0C",		-- 00dcd4: 0C10             RRC     R12
						   56533 => x"F0",
						   56534 => x"30",		-- 00dcd6: 3041             RET     
						   56535 => x"21",
						   -- Begin: __mspabi_slll_15
						   56536 => x"0C",		-- 00dcd8: 0C5C             RLA.W   R12
						   56537 => x"3C",
						   56538 => x"0D",		-- 00dcda: 0D6D             RLC.W   R13
						   56539 => x"4D",
						   -- Begin: __mspabi_slll_14
						   56540 => x"0C",		-- 00dcdc: 0C5C             RLA.W   R12
						   56541 => x"3C",
						   56542 => x"0D",		-- 00dcde: 0D6D             RLC.W   R13
						   56543 => x"4D",
						   -- Begin: __mspabi_slll_13
						   56544 => x"0C",		-- 00dce0: 0C5C             RLA.W   R12
						   56545 => x"3C",
						   56546 => x"0D",		-- 00dce2: 0D6D             RLC.W   R13
						   56547 => x"4D",
						   -- Begin: __mspabi_slll_12
						   56548 => x"0C",		-- 00dce4: 0C5C             RLA.W   R12
						   56549 => x"3C",
						   56550 => x"0D",		-- 00dce6: 0D6D             RLC.W   R13
						   56551 => x"4D",
						   -- Begin: __mspabi_slll_11
						   56552 => x"0C",		-- 00dce8: 0C5C             RLA.W   R12
						   56553 => x"3C",
						   56554 => x"0D",		-- 00dcea: 0D6D             RLC.W   R13
						   56555 => x"4D",
						   -- Begin: __mspabi_slll_10
						   56556 => x"0C",		-- 00dcec: 0C5C             RLA.W   R12
						   56557 => x"3C",
						   56558 => x"0D",		-- 00dcee: 0D6D             RLC.W   R13
						   56559 => x"4D",
						   -- Begin: __mspabi_slll_9
						   56560 => x"0C",		-- 00dcf0: 0C5C             RLA.W   R12
						   56561 => x"3C",
						   56562 => x"0D",		-- 00dcf2: 0D6D             RLC.W   R13
						   56563 => x"4D",
						   -- Begin: __mspabi_slll_8
						   56564 => x"0C",		-- 00dcf4: 0C5C             RLA.W   R12
						   56565 => x"3C",
						   56566 => x"0D",		-- 00dcf6: 0D6D             RLC.W   R13
						   56567 => x"4D",
						   -- Begin: __mspabi_slll_7
						   56568 => x"0C",		-- 00dcf8: 0C5C             RLA.W   R12
						   56569 => x"3C",
						   56570 => x"0D",		-- 00dcfa: 0D6D             RLC.W   R13
						   56571 => x"4D",
						   -- Begin: __mspabi_slll_6
						   56572 => x"0C",		-- 00dcfc: 0C5C             RLA.W   R12
						   56573 => x"3C",
						   56574 => x"0D",		-- 00dcfe: 0D6D             RLC.W   R13
						   56575 => x"4D",
						   -- Begin: __mspabi_slll_5
						   56576 => x"0C",		-- 00dd00: 0C5C             RLA.W   R12
						   56577 => x"3C",
						   56578 => x"0D",		-- 00dd02: 0D6D             RLC.W   R13
						   56579 => x"4D",
						   -- Begin: __mspabi_slll_4
						   56580 => x"0C",		-- 00dd04: 0C5C             RLA.W   R12
						   56581 => x"3C",
						   56582 => x"0D",		-- 00dd06: 0D6D             RLC.W   R13
						   56583 => x"4D",
						   -- Begin: __mspabi_slll_3
						   56584 => x"0C",		-- 00dd08: 0C5C             RLA.W   R12
						   56585 => x"3C",
						   56586 => x"0D",		-- 00dd0a: 0D6D             RLC.W   R13
						   56587 => x"4D",
						   -- Begin: __mspabi_slll_2
						   56588 => x"0C",		-- 00dd0c: 0C5C             RLA.W   R12
						   56589 => x"3C",
						   56590 => x"0D",		-- 00dd0e: 0D6D             RLC.W   R13
						   56591 => x"4D",
						   -- Begin: __mspabi_slll_1
						   56592 => x"0C",		-- 00dd10: 0C5C             RLA.W   R12
						   56593 => x"3C",
						   56594 => x"0D",		-- 00dd12: 0D6D             RLC.W   R13
						   56595 => x"4D",
						   56596 => x"30",		-- 00dd14: 3041             RET     
						   56597 => x"21",
						   -- Begin: printf
						   56598 => x"0A",		-- 00dd16: 0A12             PUSH    R10
						   56599 => x"F2",
						   56600 => x"21",		-- 00dd18: 2183             DECD.W  SP
						   56601 => x"63",
						   56602 => x"92",		-- 00dd1a: 9212             CALL    &_lock
						   56603 => x"F2",
						   56604 => x"F2",		-- 00dd1c: F220            
						   56605 => x"20",
						   56606 => x"B2",		-- 00dd1e: B293             CMP.W   #-1,&0x200c
						   56607 => x"73",
						   56608 => x"0C",		-- 00dd20: 0C20            
						   56609 => x"20",
						   56610 => x"02",		-- 00dd22: 0220             JNE     ($C$L1)
						   56611 => x"00",
						   56612 => x"3A",		-- 00dd24: 3A43             MOV.W   #-1,R10
						   56613 => x"23",
						   56614 => x"0F",		-- 00dd26: 0F3C             JMP     ($C$L2)
						   56615 => x"1C",
						   56616 => x"B1",		-- 00dd28: B140             MOV.W   #0xe1f8,0x0000(SP)
						   56617 => x"20",
						   56618 => x"F8",		-- 00dd2a: F8E1            
						   56619 => x"E1",
						   56620 => x"00",		-- 00dd2c: 0000            
						   56621 => x"00",
						   56622 => x"0D",		-- 00dd2e: 0D41             MOV.W   SP,R13
						   56623 => x"21",
						   56624 => x"3D",		-- 00dd30: 3D52             ADD.W   #8,R13
						   56625 => x"32",
						   56626 => x"3E",		-- 00dd32: 3E40             MOV.W   #0x200c,R14
						   56627 => x"20",
						   56628 => x"0C",		-- 00dd34: 0C20            
						   56629 => x"20",
						   56630 => x"0C",		-- 00dd36: 0C41             MOV.W   SP,R12
						   56631 => x"21",
						   56632 => x"3C",		-- 00dd38: 3C50             ADD.W   #0x0006,R12
						   56633 => x"30",
						   56634 => x"06",		-- 00dd3a: 0600            
						   56635 => x"00",
						   56636 => x"3F",		-- 00dd3c: 3F40             MOV.W   #0xe1ec,R15
						   56637 => x"20",
						   56638 => x"EC",		-- 00dd3e: ECE1            
						   56639 => x"E1",
						   56640 => x"B0",		-- 00dd40: B012             CALL    #__TI_printfi
						   56641 => x"F2",
						   56642 => x"2C",		-- 00dd42: 2CAC            
						   56643 => x"AC",
						   56644 => x"0A",		-- 00dd44: 0A4C             MOV.W   R12,R10
						   56645 => x"2C",
						   56646 => x"92",		-- 00dd46: 9212             CALL    &_unlock
						   56647 => x"F2",
						   56648 => x"F4",		-- 00dd48: F420            
						   56649 => x"20",
						   56650 => x"0C",		-- 00dd4a: 0C4A             MOV.W   R10,R12
						   56651 => x"2A",
						   56652 => x"21",		-- 00dd4c: 2153             INCD.W  SP
						   56653 => x"33",
						   56654 => x"3A",		-- 00dd4e: 3A41             POP.W   R10
						   56655 => x"21",
						   56656 => x"30",		-- 00dd50: 3041             RET     
						   56657 => x"21",
						   -- Begin: __TI_cleanup
						   56658 => x"0A",		-- 00dd52: 0A12             PUSH    R10
						   56659 => x"F2",
						   56660 => x"09",		-- 00dd54: 0912             PUSH    R9
						   56661 => x"F2",
						   56662 => x"3C",		-- 00dd56: 3C40             MOV.W   #0x2000,R12
						   56663 => x"20",
						   56664 => x"00",		-- 00dd58: 0020            
						   56665 => x"20",
						   56666 => x"B0",		-- 00dd5a: B012             CALL    #__TI_closefile
						   56667 => x"F2",
						   56668 => x"30",		-- 00dd5c: 30D4            
						   56669 => x"D4",
						   56670 => x"A2",		-- 00dd5e: A293             CMP.W   #2,&__TI_ft_end
						   56671 => x"73",
						   56672 => x"F6",		-- 00dd60: F620            
						   56673 => x"20",
						   56674 => x"0F",		-- 00dd62: 0F38             JL      ($C$L37)
						   56675 => x"18",
						   56676 => x"3A",		-- 00dd64: 3A40             MOV.W   #0x200c,R10
						   56677 => x"20",
						   56678 => x"0C",		-- 00dd66: 0C20            
						   56679 => x"20",
						   56680 => x"19",		-- 00dd68: 1943             MOV.W   #1,R9
						   56681 => x"23",
						   56682 => x"8A",		-- 00dd6a: 8A93             TST.W   0x0000(R10)
						   56683 => x"73",
						   56684 => x"00",		-- 00dd6c: 0000            
						   56685 => x"00",
						   56686 => x"03",		-- 00dd6e: 0338             JL      ($C$L36)
						   56687 => x"18",
						   56688 => x"0C",		-- 00dd70: 0C4A             MOV.W   R10,R12
						   56689 => x"2A",
						   56690 => x"B0",		-- 00dd72: B012             CALL    #__TI_closefile
						   56691 => x"F2",
						   56692 => x"30",		-- 00dd74: 30D4            
						   56693 => x"D4",
						   56694 => x"3A",		-- 00dd76: 3A50             ADD.W   #0x000c,R10
						   56695 => x"30",
						   56696 => x"0C",		-- 00dd78: 0C00            
						   56697 => x"00",
						   56698 => x"19",		-- 00dd7a: 1953             INC.W   R9
						   56699 => x"33",
						   56700 => x"19",		-- 00dd7c: 1992             CMP.W   &__TI_ft_end,R9
						   56701 => x"72",
						   56702 => x"F6",		-- 00dd7e: F620            
						   56703 => x"20",
						   56704 => x"F4",		-- 00dd80: F43B             JL      ($C$L35)
						   56705 => x"1B",
						   56706 => x"30",		-- 00dd82: 3040             BR      #__mspabi_func_epilog_2
						   56707 => x"20",
						   56708 => x"9E",		-- 00dd84: 9EE1            
						   56709 => x"E1",
						   -- Begin: finddevice
						   56710 => x"0A",		-- 00dd86: 0A12             PUSH    R10
						   56711 => x"F2",
						   56712 => x"09",		-- 00dd88: 0912             PUSH    R9
						   56713 => x"F2",
						   56714 => x"08",		-- 00dd8a: 0812             PUSH    R8
						   56715 => x"F2",
						   56716 => x"08",		-- 00dd8c: 084C             MOV.W   R12,R8
						   56717 => x"2C",
						   56718 => x"C8",		-- 00dd8e: C893             TST.B   0x0000(R8)
						   56719 => x"73",
						   56720 => x"00",		-- 00dd90: 0000            
						   56721 => x"00",
						   56722 => x"10",		-- 00dd92: 1024             JEQ     ($C$L3)
						   56723 => x"04",
						   56724 => x"3A",		-- 00dd94: 3A40             MOV.W   #0x2092,R10
						   56725 => x"20",
						   56726 => x"92",		-- 00dd96: 9220            
						   56727 => x"20",
						   56728 => x"29",		-- 00dd98: 2943             MOV.W   #2,R9
						   56729 => x"23",
						   56730 => x"0C",		-- 00dd9a: 0C4A             MOV.W   R10,R12
						   56731 => x"2A",
						   56732 => x"0D",		-- 00dd9c: 0D48             MOV.W   R8,R13
						   56733 => x"28",
						   56734 => x"B0",		-- 00dd9e: B012             CALL    #strcmp
						   56735 => x"F2",
						   56736 => x"BA",		-- 00dda0: BAE0            
						   56737 => x"E0",
						   56738 => x"0C",		-- 00dda2: 0C93             TST.W   R12
						   56739 => x"73",
						   56740 => x"03",		-- 00dda4: 0320             JNE     ($C$L2)
						   56741 => x"00",
						   56742 => x"0C",		-- 00dda6: 0C4A             MOV.W   R10,R12
						   56743 => x"2A",
						   56744 => x"30",		-- 00dda8: 3040             BR      #__mspabi_func_epilog_3
						   56745 => x"20",
						   56746 => x"9C",		-- 00ddaa: 9CE1            
						   56747 => x"E1",
						   56748 => x"3A",		-- 00ddac: 3A50             ADD.W   #0x001a,R10
						   56749 => x"30",
						   56750 => x"1A",		-- 00ddae: 1A00            
						   56751 => x"00",
						   56752 => x"19",		-- 00ddb0: 1983             DEC.W   R9
						   56753 => x"63",
						   56754 => x"F3",		-- 00ddb2: F323             JNE     ($C$L1)
						   56755 => x"03",
						   56756 => x"0C",		-- 00ddb4: 0C43             CLR.W   R12
						   56757 => x"23",
						   56758 => x"30",		-- 00ddb6: 3040             BR      #__mspabi_func_epilog_3
						   56759 => x"20",
						   56760 => x"9C",		-- 00ddb8: 9CE1            
						   56761 => x"E1",
						   -- Begin: __TI_writemsg
						   56762 => x"82",		-- 00ddba: 824F             MOV.W   R15,&_CIOBUF_
						   56763 => x"2F",
						   56764 => x"00",		-- 00ddbc: 0080            
						   56765 => x"80",
						   56766 => x"C2",		-- 00ddbe: C24C             MOV.B   R12,&0x8002
						   56767 => x"2C",
						   56768 => x"02",		-- 00ddc0: 0280            
						   56769 => x"80",
						   56770 => x"3C",		-- 00ddc2: 3C40             MOV.W   #0x8003,R12
						   56771 => x"20",
						   56772 => x"03",		-- 00ddc4: 0380            
						   56773 => x"80",
						   56774 => x"3B",		-- 00ddc6: 3B42             MOV.W   #8,R11
						   56775 => x"22",
						   56776 => x"1C",		-- 00ddc8: 1C53             INC.W   R12
						   56777 => x"33",
						   56778 => x"FC",		-- 00ddca: FC4D             MOV.B   @R13+,0xffff(R12)
						   56779 => x"2D",
						   56780 => x"FF",		-- 00ddcc: FFFF            
						   56781 => x"FF",
						   56782 => x"1B",		-- 00ddce: 1B83             DEC.W   R11
						   56783 => x"63",
						   56784 => x"FB",		-- 00ddd0: FB23             JNE     ($C$L1)
						   56785 => x"03",
						   56786 => x"0F",		-- 00ddd2: 0F93             TST.W   R15
						   56787 => x"73",
						   56788 => x"07",		-- 00ddd4: 0724             JEQ     (C$$IO$$)
						   56789 => x"04",
						   56790 => x"3D",		-- 00ddd6: 3D40             MOV.W   #0x800b,R13
						   56791 => x"20",
						   56792 => x"0B",		-- 00ddd8: 0B80            
						   56793 => x"80",
						   56794 => x"1D",		-- 00ddda: 1D53             INC.W   R13
						   56795 => x"33",
						   56796 => x"FD",		-- 00dddc: FD4E             MOV.B   @R14+,0xffff(R13)
						   56797 => x"2E",
						   56798 => x"FF",		-- 00ddde: FFFF            
						   56799 => x"FF",
						   56800 => x"1F",		-- 00dde0: 1F83             DEC.W   R15
						   56801 => x"63",
						   56802 => x"FB",		-- 00dde2: FB23             JNE     ($C$L2)
						   56803 => x"03",
						   56804 => x"03",		-- 00dde4: 0343             NOP     
						   56805 => x"23",
						   56806 => x"30",		-- 00dde6: 3041             RET     
						   56807 => x"21",
						   -- Begin: __mspabi_subd
						   56808 => x"31",		-- 00dde8: 3182             SUB.W   #8,SP
						   56809 => x"62",
						   56810 => x"81",		-- 00ddea: 814C             MOV.W   R12,0x0000(SP)
						   56811 => x"2C",
						   56812 => x"00",		-- 00ddec: 0000            
						   56813 => x"00",
						   56814 => x"81",		-- 00ddee: 814D             MOV.W   R13,0x0002(SP)
						   56815 => x"2D",
						   56816 => x"02",		-- 00ddf0: 0200            
						   56817 => x"00",
						   56818 => x"81",		-- 00ddf2: 814E             MOV.W   R14,0x0004(SP)
						   56819 => x"2E",
						   56820 => x"04",		-- 00ddf4: 0400            
						   56821 => x"00",
						   56822 => x"81",		-- 00ddf6: 814F             MOV.W   R15,0x0006(SP)
						   56823 => x"2F",
						   56824 => x"06",		-- 00ddf8: 0600            
						   56825 => x"00",
						   56826 => x"F1",		-- 00ddfa: F1E0             XOR.B   #0x0080,0x0007(SP)
						   56827 => x"C0",
						   56828 => x"80",		-- 00ddfc: 8000            
						   56829 => x"00",
						   56830 => x"07",		-- 00ddfe: 0700            
						   56831 => x"00",
						   56832 => x"2C",		-- 00de00: 2C41             MOV.W   @SP,R12
						   56833 => x"21",
						   56834 => x"1D",		-- 00de02: 1D41             MOV.W   0x0002(SP),R13
						   56835 => x"21",
						   56836 => x"02",		-- 00de04: 0200            
						   56837 => x"00",
						   56838 => x"1E",		-- 00de06: 1E41             MOV.W   0x0004(SP),R14
						   56839 => x"21",
						   56840 => x"04",		-- 00de08: 0400            
						   56841 => x"00",
						   56842 => x"1F",		-- 00de0a: 1F41             MOV.W   0x0006(SP),R15
						   56843 => x"21",
						   56844 => x"06",		-- 00de0c: 0600            
						   56845 => x"00",
						   56846 => x"B0",		-- 00de0e: B012             CALL    #__mspabi_addd
						   56847 => x"F2",
						   56848 => x"5E",		-- 00de10: 5E9A            
						   56849 => x"9A",
						   56850 => x"31",		-- 00de12: 3152             ADD.W   #8,SP
						   56851 => x"32",
						   56852 => x"30",		-- 00de14: 3041             RET     
						   56853 => x"21",
						   -- Begin: copysignl
						   -- Begin: copysign
						   56854 => x"0A",		-- 00de16: 0A12             PUSH    R10
						   56855 => x"F2",
						   56856 => x"1A",		-- 00de18: 1A41             MOV.W   0x0008(SP),R10
						   56857 => x"21",
						   56858 => x"08",		-- 00de1a: 0800            
						   56859 => x"00",
						   56860 => x"1B",		-- 00de1c: 1B41             MOV.W   0x000a(SP),R11
						   56861 => x"21",
						   56862 => x"0A",		-- 00de1e: 0A00            
						   56863 => x"00",
						   56864 => x"0A",		-- 00de20: 0AF3             AND.W   #0,R10
						   56865 => x"D3",
						   56866 => x"3B",		-- 00de22: 3BF0             AND.W   #0x8000,R11
						   56867 => x"D0",
						   56868 => x"00",		-- 00de24: 0080            
						   56869 => x"80",
						   56870 => x"3E",		-- 00de26: 3EF3             AND.W   #-1,R14
						   56871 => x"D3",
						   56872 => x"3F",		-- 00de28: 3FF0             AND.W   #0x7fff,R15
						   56873 => x"D0",
						   56874 => x"FF",		-- 00de2a: FF7F            
						   56875 => x"7F",
						   56876 => x"0E",		-- 00de2c: 0EDA             BIS.W   R10,R14
						   56877 => x"BA",
						   56878 => x"0F",		-- 00de2e: 0FDB             BIS.W   R11,R15
						   56879 => x"BB",
						   56880 => x"0B",		-- 00de30: 0B43             CLR.W   R11
						   56881 => x"23",
						   56882 => x"0B",		-- 00de32: 0BDD             BIS.W   R13,R11
						   56883 => x"BD",
						   56884 => x"0D",		-- 00de34: 0D43             CLR.W   R13
						   56885 => x"23",
						   56886 => x"0D",		-- 00de36: 0DDC             BIS.W   R12,R13
						   56887 => x"BC",
						   56888 => x"0E",		-- 00de38: 0ED3             BIS.W   #0,R14
						   56889 => x"B3",
						   56890 => x"0F",		-- 00de3a: 0FD3             BIS.W   #0,R15
						   56891 => x"B3",
						   56892 => x"0C",		-- 00de3c: 0C4D             MOV.W   R13,R12
						   56893 => x"2D",
						   56894 => x"0D",		-- 00de3e: 0D4B             MOV.W   R11,R13
						   56895 => x"2B",
						   56896 => x"3A",		-- 00de40: 3A41             POP.W   R10
						   56897 => x"21",
						   56898 => x"30",		-- 00de42: 3041             RET     
						   56899 => x"21",
						   -- Begin: __TI_readmsg
						   56900 => x"1F",		-- 00de44: 1F42             MOV.W   &_CIOBUF_,R15
						   56901 => x"22",
						   56902 => x"00",		-- 00de46: 0080            
						   56903 => x"80",
						   56904 => x"3B",		-- 00de48: 3B40             MOV.W   #0x8002,R11
						   56905 => x"20",
						   56906 => x"02",		-- 00de4a: 0280            
						   56907 => x"80",
						   56908 => x"3E",		-- 00de4c: 3E42             MOV.W   #8,R14
						   56909 => x"22",
						   56910 => x"1C",		-- 00de4e: 1C53             INC.W   R12
						   56911 => x"33",
						   56912 => x"FC",		-- 00de50: FC4B             MOV.B   @R11+,0xffff(R12)
						   56913 => x"2B",
						   56914 => x"FF",		-- 00de52: FFFF            
						   56915 => x"FF",
						   56916 => x"1E",		-- 00de54: 1E83             DEC.W   R14
						   56917 => x"63",
						   56918 => x"FB",		-- 00de56: FB23             JNE     ($C$L4)
						   56919 => x"03",
						   56920 => x"0D",		-- 00de58: 0D93             TST.W   R13
						   56921 => x"73",
						   56922 => x"09",		-- 00de5a: 0924             JEQ     ($C$L6)
						   56923 => x"04",
						   56924 => x"0F",		-- 00de5c: 0F93             TST.W   R15
						   56925 => x"73",
						   56926 => x"07",		-- 00de5e: 0724             JEQ     ($C$L6)
						   56927 => x"04",
						   56928 => x"3E",		-- 00de60: 3E40             MOV.W   #0x800a,R14
						   56929 => x"20",
						   56930 => x"0A",		-- 00de62: 0A80            
						   56931 => x"80",
						   56932 => x"1D",		-- 00de64: 1D53             INC.W   R13
						   56933 => x"33",
						   56934 => x"FD",		-- 00de66: FD4E             MOV.B   @R14+,0xffff(R13)
						   56935 => x"2E",
						   56936 => x"FF",		-- 00de68: FFFF            
						   56937 => x"FF",
						   56938 => x"1F",		-- 00de6a: 1F83             DEC.W   R15
						   56939 => x"63",
						   56940 => x"FB",		-- 00de6c: FB23             JNE     ($C$L5)
						   56941 => x"03",
						   56942 => x"30",		-- 00de6e: 3041             RET     
						   56943 => x"21",
						   -- Begin: __mspabi_srai
						   56944 => x"3D",		-- 00de70: 3DF0             AND.W   #0x000f,R13
						   56945 => x"D0",
						   56946 => x"0F",		-- 00de72: 0F00            
						   56947 => x"00",
						   56948 => x"3D",		-- 00de74: 3DE0             XOR.W   #0x000f,R13
						   56949 => x"C0",
						   56950 => x"0F",		-- 00de76: 0F00            
						   56951 => x"00",
						   56952 => x"0D",		-- 00de78: 0D5D             RLA.W   R13
						   56953 => x"3D",
						   56954 => x"00",		-- 00de7a: 005D             ADD.W   R13,PC
						   56955 => x"3D",
						   -- Begin: __mspabi_srai_15
						   56956 => x"0C",		-- 00de7c: 0C11             RRA     R12
						   56957 => x"F1",
						   -- Begin: __mspabi_srai_14
						   56958 => x"0C",		-- 00de7e: 0C11             RRA     R12
						   56959 => x"F1",
						   -- Begin: __mspabi_srai_13
						   56960 => x"0C",		-- 00de80: 0C11             RRA     R12
						   56961 => x"F1",
						   -- Begin: __mspabi_srai_12
						   56962 => x"0C",		-- 00de82: 0C11             RRA     R12
						   56963 => x"F1",
						   -- Begin: __mspabi_srai_11
						   56964 => x"0C",		-- 00de84: 0C11             RRA     R12
						   56965 => x"F1",
						   -- Begin: __mspabi_srai_10
						   56966 => x"0C",		-- 00de86: 0C11             RRA     R12
						   56967 => x"F1",
						   -- Begin: __mspabi_srai_9
						   56968 => x"0C",		-- 00de88: 0C11             RRA     R12
						   56969 => x"F1",
						   -- Begin: __mspabi_srai_8
						   56970 => x"0C",		-- 00de8a: 0C11             RRA     R12
						   56971 => x"F1",
						   -- Begin: __mspabi_srai_7
						   56972 => x"0C",		-- 00de8c: 0C11             RRA     R12
						   56973 => x"F1",
						   -- Begin: __mspabi_srai_6
						   56974 => x"0C",		-- 00de8e: 0C11             RRA     R12
						   56975 => x"F1",
						   -- Begin: __mspabi_srai_5
						   56976 => x"0C",		-- 00de90: 0C11             RRA     R12
						   56977 => x"F1",
						   -- Begin: __mspabi_srai_4
						   56978 => x"0C",		-- 00de92: 0C11             RRA     R12
						   56979 => x"F1",
						   -- Begin: __mspabi_srai_3
						   56980 => x"0C",		-- 00de94: 0C11             RRA     R12
						   56981 => x"F1",
						   -- Begin: __mspabi_srai_2
						   56982 => x"0C",		-- 00de96: 0C11             RRA     R12
						   56983 => x"F1",
						   -- Begin: __mspabi_srai_1
						   56984 => x"0C",		-- 00de98: 0C11             RRA     R12
						   56985 => x"F1",
						   56986 => x"30",		-- 00de9a: 3041             RET     
						   56987 => x"21",
						   -- Begin: __mspabi_slli
						   56988 => x"3D",		-- 00de9c: 3DF0             AND.W   #0x000f,R13
						   56989 => x"D0",
						   56990 => x"0F",		-- 00de9e: 0F00            
						   56991 => x"00",
						   56992 => x"3D",		-- 00dea0: 3DE0             XOR.W   #0x000f,R13
						   56993 => x"C0",
						   56994 => x"0F",		-- 00dea2: 0F00            
						   56995 => x"00",
						   56996 => x"0D",		-- 00dea4: 0D5D             RLA.W   R13
						   56997 => x"3D",
						   56998 => x"00",		-- 00dea6: 005D             ADD.W   R13,PC
						   56999 => x"3D",
						   -- Begin: __mspabi_slli_15
						   57000 => x"0C",		-- 00dea8: 0C5C             RLA.W   R12
						   57001 => x"3C",
						   -- Begin: __mspabi_slli_14
						   57002 => x"0C",		-- 00deaa: 0C5C             RLA.W   R12
						   57003 => x"3C",
						   -- Begin: __mspabi_slli_13
						   57004 => x"0C",		-- 00deac: 0C5C             RLA.W   R12
						   57005 => x"3C",
						   -- Begin: __mspabi_slli_12
						   57006 => x"0C",		-- 00deae: 0C5C             RLA.W   R12
						   57007 => x"3C",
						   -- Begin: __mspabi_slli_11
						   57008 => x"0C",		-- 00deb0: 0C5C             RLA.W   R12
						   57009 => x"3C",
						   -- Begin: __mspabi_slli_10
						   57010 => x"0C",		-- 00deb2: 0C5C             RLA.W   R12
						   57011 => x"3C",
						   -- Begin: __mspabi_slli_9
						   57012 => x"0C",		-- 00deb4: 0C5C             RLA.W   R12
						   57013 => x"3C",
						   -- Begin: __mspabi_slli_8
						   57014 => x"0C",		-- 00deb6: 0C5C             RLA.W   R12
						   57015 => x"3C",
						   -- Begin: __mspabi_slli_7
						   57016 => x"0C",		-- 00deb8: 0C5C             RLA.W   R12
						   57017 => x"3C",
						   -- Begin: __mspabi_slli_6
						   57018 => x"0C",		-- 00deba: 0C5C             RLA.W   R12
						   57019 => x"3C",
						   -- Begin: __mspabi_slli_5
						   57020 => x"0C",		-- 00debc: 0C5C             RLA.W   R12
						   57021 => x"3C",
						   -- Begin: __mspabi_slli_4
						   57022 => x"0C",		-- 00debe: 0C5C             RLA.W   R12
						   57023 => x"3C",
						   -- Begin: __mspabi_slli_3
						   57024 => x"0C",		-- 00dec0: 0C5C             RLA.W   R12
						   57025 => x"3C",
						   -- Begin: __mspabi_slli_2
						   57026 => x"0C",		-- 00dec2: 0C5C             RLA.W   R12
						   57027 => x"3C",
						   -- Begin: __mspabi_slli_1
						   57028 => x"0C",		-- 00dec4: 0C5C             RLA.W   R12
						   57029 => x"3C",
						   57030 => x"30",		-- 00dec6: 3041             RET     
						   57031 => x"21",
						   -- Begin: strncpy
						   57032 => x"0E",		-- 00dec8: 0E93             TST.W   R14
						   57033 => x"73",
						   57034 => x"13",		-- 00deca: 1324             JEQ     ($C$L4)
						   57035 => x"04",
						   57036 => x"0F",		-- 00decc: 0F4C             MOV.W   R12,R15
						   57037 => x"2C",
						   57038 => x"6B",		-- 00dece: 6B4D             MOV.B   @R13,R11
						   57039 => x"2D",
						   57040 => x"1F",		-- 00ded0: 1F53             INC.W   R15
						   57041 => x"33",
						   57042 => x"CF",		-- 00ded2: CF4B             MOV.B   R11,0xffff(R15)
						   57043 => x"2B",
						   57044 => x"FF",		-- 00ded4: FFFF            
						   57045 => x"FF",
						   57046 => x"0B",		-- 00ded6: 0B93             TST.W   R11
						   57047 => x"73",
						   57048 => x"03",		-- 00ded8: 0324             JEQ     ($C$L2)
						   57049 => x"04",
						   57050 => x"1D",		-- 00deda: 1D53             INC.W   R13
						   57051 => x"33",
						   57052 => x"1E",		-- 00dedc: 1E83             DEC.W   R14
						   57053 => x"63",
						   57054 => x"F7",		-- 00dede: F723             JNE     ($C$L1)
						   57055 => x"03",
						   57056 => x"0D",		-- 00dee0: 0D4E             MOV.W   R14,R13
						   57057 => x"2E",
						   57058 => x"1E",		-- 00dee2: 1E83             DEC.W   R14
						   57059 => x"63",
						   57060 => x"2D",		-- 00dee4: 2D93             CMP.W   #2,R13
						   57061 => x"73",
						   57062 => x"05",		-- 00dee6: 0528             JLO     ($C$L4)
						   57063 => x"08",
						   57064 => x"1F",		-- 00dee8: 1F53             INC.W   R15
						   57065 => x"33",
						   57066 => x"CF",		-- 00deea: CF43             CLR.B   0xffff(R15)
						   57067 => x"23",
						   57068 => x"FF",		-- 00deec: FFFF            
						   57069 => x"FF",
						   57070 => x"1E",		-- 00deee: 1E83             DEC.W   R14
						   57071 => x"63",
						   57072 => x"FB",		-- 00def0: FB23             JNE     ($C$L3)
						   57073 => x"03",
						   57074 => x"30",		-- 00def2: 3041             RET     
						   57075 => x"21",
						   -- Begin: __mspabi_negd
						   57076 => x"31",		-- 00def4: 3182             SUB.W   #8,SP
						   57077 => x"62",
						   57078 => x"81",		-- 00def6: 814C             MOV.W   R12,0x0000(SP)
						   57079 => x"2C",
						   57080 => x"00",		-- 00def8: 0000            
						   57081 => x"00",
						   57082 => x"81",		-- 00defa: 814D             MOV.W   R13,0x0002(SP)
						   57083 => x"2D",
						   57084 => x"02",		-- 00defc: 0200            
						   57085 => x"00",
						   57086 => x"81",		-- 00defe: 814E             MOV.W   R14,0x0004(SP)
						   57087 => x"2E",
						   57088 => x"04",		-- 00df00: 0400            
						   57089 => x"00",
						   57090 => x"81",		-- 00df02: 814F             MOV.W   R15,0x0006(SP)
						   57091 => x"2F",
						   57092 => x"06",		-- 00df04: 0600            
						   57093 => x"00",
						   57094 => x"F1",		-- 00df06: F1E0             XOR.B   #0x0080,0x0007(SP)
						   57095 => x"C0",
						   57096 => x"80",		-- 00df08: 8000            
						   57097 => x"00",
						   57098 => x"07",		-- 00df0a: 0700            
						   57099 => x"00",
						   57100 => x"2C",		-- 00df0c: 2C41             MOV.W   @SP,R12
						   57101 => x"21",
						   57102 => x"1D",		-- 00df0e: 1D41             MOV.W   0x0002(SP),R13
						   57103 => x"21",
						   57104 => x"02",		-- 00df10: 0200            
						   57105 => x"00",
						   57106 => x"1E",		-- 00df12: 1E41             MOV.W   0x0004(SP),R14
						   57107 => x"21",
						   57108 => x"04",		-- 00df14: 0400            
						   57109 => x"00",
						   57110 => x"1F",		-- 00df16: 1F41             MOV.W   0x0006(SP),R15
						   57111 => x"21",
						   57112 => x"06",		-- 00df18: 0600            
						   57113 => x"00",
						   57114 => x"31",		-- 00df1a: 3152             ADD.W   #8,SP
						   57115 => x"32",
						   57116 => x"30",		-- 00df1c: 3041             RET     
						   57117 => x"21",
						   -- Begin: __mspabi_fixdi
						   57118 => x"B0",		-- 00df1e: B012             CALL    #__mspabi_fixdli
						   57119 => x"F2",
						   57120 => x"A2",		-- 00df20: A2D4            
						   57121 => x"D4",
						   57122 => x"0D",		-- 00df22: 0D93             TST.W   R13
						   57123 => x"73",
						   57124 => x"07",		-- 00df24: 0738             JL      ($C$L7)
						   57125 => x"18",
						   57126 => x"03",		-- 00df26: 0320             JNE     ($C$L6)
						   57127 => x"00",
						   57128 => x"3C",		-- 00df28: 3C90             CMP.W   #0x8000,R12
						   57129 => x"70",
						   57130 => x"00",		-- 00df2a: 0080            
						   57131 => x"80",
						   57132 => x"03",		-- 00df2c: 0328             JLO     ($C$L7)
						   57133 => x"08",
						   57134 => x"3C",		-- 00df2e: 3C40             MOV.W   #0x7fff,R12
						   57135 => x"20",
						   57136 => x"FF",		-- 00df30: FF7F            
						   57137 => x"7F",
						   57138 => x"30",		-- 00df32: 3041             RET     
						   57139 => x"21",
						   57140 => x"3D",		-- 00df34: 3D93             CMP.W   #-1,R13
						   57141 => x"73",
						   57142 => x"04",		-- 00df36: 0438             JL      ($C$L8)
						   57143 => x"18",
						   57144 => x"05",		-- 00df38: 0520             JNE     ($C$L9)
						   57145 => x"00",
						   57146 => x"3C",		-- 00df3a: 3C90             CMP.W   #0x8000,R12
						   57147 => x"70",
						   57148 => x"00",		-- 00df3c: 0080            
						   57149 => x"80",
						   57150 => x"02",		-- 00df3e: 022C             JHS     ($C$L9)
						   57151 => x"0C",
						   57152 => x"3C",		-- 00df40: 3C40             MOV.W   #0x8000,R12
						   57153 => x"20",
						   57154 => x"00",		-- 00df42: 0080            
						   57155 => x"80",
						   57156 => x"30",		-- 00df44: 3041             RET     
						   57157 => x"21",
						   -- Begin: free_list_insert
						   57158 => x"2F",		-- 00df46: 2F4C             MOV.W   @R12,R15
						   57159 => x"2C",
						   57160 => x"1F",		-- 00df48: 1FC3             BIC.W   #1,R15
						   57161 => x"A3",
						   57162 => x"3E",		-- 00df4a: 3E40             MOV.W   #0x21a6,R14
						   57163 => x"20",
						   57164 => x"A6",		-- 00df4c: A621            
						   57165 => x"21",
						   57166 => x"03",		-- 00df4e: 033C             JMP     ($C$L5)
						   57167 => x"1C",
						   57168 => x"2D",		-- 00df50: 2D42             MOV.W   #4,R13
						   57169 => x"22",
						   57170 => x"2D",		-- 00df52: 2D5E             ADD.W   @R14,R13
						   57171 => x"3E",
						   57172 => x"0E",		-- 00df54: 0E4D             MOV.W   R13,R14
						   57173 => x"2D",
						   57174 => x"2D",		-- 00df56: 2D4E             MOV.W   @R14,R13
						   57175 => x"2E",
						   57176 => x"0D",		-- 00df58: 0D93             TST.W   R13
						   57177 => x"73",
						   57178 => x"04",		-- 00df5a: 0424             JEQ     ($C$L6)
						   57179 => x"04",
						   57180 => x"2D",		-- 00df5c: 2D4D             MOV.W   @R13,R13
						   57181 => x"2D",
						   57182 => x"1D",		-- 00df5e: 1DC3             BIC.W   #1,R13
						   57183 => x"A3",
						   57184 => x"0D",		-- 00df60: 0D9F             CMP.W   R15,R13
						   57185 => x"7F",
						   57186 => x"F6",		-- 00df62: F62B             JLO     ($C$L4)
						   57187 => x"0B",
						   57188 => x"AC",		-- 00df64: AC4E             MOV.W   @R14,0x0004(R12)
						   57189 => x"2E",
						   57190 => x"04",		-- 00df66: 0400            
						   57191 => x"00",
						   57192 => x"8E",		-- 00df68: 8E4C             MOV.W   R12,0x0000(R14)
						   57193 => x"2C",
						   57194 => x"00",		-- 00df6a: 0000            
						   57195 => x"00",
						   57196 => x"30",		-- 00df6c: 3041             RET     
						   57197 => x"21",
						   -- Begin: remove
						   -- Begin: unlink
						   57198 => x"0A",		-- 00df6e: 0A12             PUSH    R10
						   57199 => x"F2",
						   57200 => x"21",		-- 00df70: 2183             DECD.W  SP
						   57201 => x"63",
						   57202 => x"81",		-- 00df72: 814C             MOV.W   R12,0x0000(SP)
						   57203 => x"2C",
						   57204 => x"00",		-- 00df74: 0000            
						   57205 => x"00",
						   57206 => x"92",		-- 00df76: 9212             CALL    &_lock
						   57207 => x"F2",
						   57208 => x"F2",		-- 00df78: F220            
						   57209 => x"20",
						   57210 => x"0C",		-- 00df7a: 0C41             MOV.W   SP,R12
						   57211 => x"21",
						   57212 => x"B0",		-- 00df7c: B012             CALL    #getdevice
						   57213 => x"F2",
						   57214 => x"96",		-- 00df7e: 96D8            
						   57215 => x"D8",
						   57216 => x"0F",		-- 00df80: 0F4C             MOV.W   R12,R15
						   57217 => x"2C",
						   57218 => x"2C",		-- 00df82: 2C41             MOV.W   @SP,R12
						   57219 => x"21",
						   57220 => x"9F",		-- 00df84: 9F12             CALL    0x0016(R15)
						   57221 => x"F2",
						   57222 => x"16",		-- 00df86: 1600            
						   57223 => x"00",
						   57224 => x"0A",		-- 00df88: 0A4C             MOV.W   R12,R10
						   57225 => x"2C",
						   57226 => x"92",		-- 00df8a: 9212             CALL    &_unlock
						   57227 => x"F2",
						   57228 => x"F4",		-- 00df8c: F420            
						   57229 => x"20",
						   57230 => x"0C",		-- 00df8e: 0C4A             MOV.W   R10,R12
						   57231 => x"2A",
						   57232 => x"21",		-- 00df90: 2153             INCD.W  SP
						   57233 => x"33",
						   57234 => x"3A",		-- 00df92: 3A41             POP.W   R10
						   57235 => x"21",
						   57236 => x"30",		-- 00df94: 3041             RET     
						   57237 => x"21",
						   -- Begin: lseek
						   57238 => x"0C",		-- 00df96: 0C93             TST.W   R12
						   57239 => x"73",
						   57240 => x"0E",		-- 00df98: 0E38             JL      ($C$L1)
						   57241 => x"18",
						   57242 => x"3C",		-- 00df9a: 3C90             CMP.W   #0x000a,R12
						   57243 => x"70",
						   57244 => x"0A",		-- 00df9c: 0A00            
						   57245 => x"00",
						   57246 => x"0B",		-- 00df9e: 0B34             JGE     ($C$L1)
						   57247 => x"14",
						   57248 => x"0C",		-- 00dfa0: 0C5C             RLA.W   R12
						   57249 => x"3C",
						   57250 => x"0C",		-- 00dfa2: 0C5C             RLA.W   R12
						   57251 => x"3C",
						   57252 => x"3C",		-- 00dfa4: 3C50             ADD.W   #0x20c6,R12
						   57253 => x"30",
						   57254 => x"C6",		-- 00dfa6: C620            
						   57255 => x"20",
						   57256 => x"2B",		-- 00dfa8: 2B4C             MOV.W   @R12,R11
						   57257 => x"2C",
						   57258 => x"0B",		-- 00dfaa: 0B93             TST.W   R11
						   57259 => x"73",
						   57260 => x"04",		-- 00dfac: 0424             JEQ     ($C$L1)
						   57261 => x"04",
						   57262 => x"1C",		-- 00dfae: 1C4C             MOV.W   0x0002(R12),R12
						   57263 => x"2C",
						   57264 => x"02",		-- 00dfb0: 0200            
						   57265 => x"00",
						   57266 => x"10",		-- 00dfb2: 104B             BR      0x0014(R11)
						   57267 => x"2B",
						   57268 => x"14",		-- 00dfb4: 1400            
						   57269 => x"00",
						   57270 => x"3C",		-- 00dfb6: 3C43             MOV.W   #-1,R12
						   57271 => x"23",
						   57272 => x"3D",		-- 00dfb8: 3D43             MOV.W   #-1,R13
						   57273 => x"23",
						   57274 => x"30",		-- 00dfba: 3041             RET     
						   57275 => x"21",
						   -- Begin: __mspabi_mpyl
						   -- Begin: __mspabi_mpyl_sw
						   57276 => x"0A",		-- 00dfbc: 0A12             PUSH    R10
						   57277 => x"F2",
						   57278 => x"0A",		-- 00dfbe: 0A43             CLR.W   R10
						   57279 => x"23",
						   57280 => x"0B",		-- 00dfc0: 0B43             CLR.W   R11
						   57281 => x"23",
						   -- Begin: mpyl_add_loop
						   57282 => x"12",		-- 00dfc2: 12C3             CLRC    
						   57283 => x"A3",
						   57284 => x"0D",		-- 00dfc4: 0D10             RRC     R13
						   57285 => x"F0",
						   57286 => x"0C",		-- 00dfc6: 0C10             RRC     R12
						   57287 => x"F0",
						   57288 => x"02",		-- 00dfc8: 0228             JLO     (shift_test_mpyl)
						   57289 => x"08",
						   57290 => x"0A",		-- 00dfca: 0A5E             ADD.W   R14,R10
						   57291 => x"3E",
						   57292 => x"0B",		-- 00dfcc: 0B6F             ADDC.W  R15,R11
						   57293 => x"4F",
						   -- Begin: shift_test_mpyl
						   57294 => x"0E",		-- 00dfce: 0E5E             RLA.W   R14
						   57295 => x"3E",
						   57296 => x"0F",		-- 00dfd0: 0F6F             RLC.W   R15
						   57297 => x"4F",
						   57298 => x"0D",		-- 00dfd2: 0D93             TST.W   R13
						   57299 => x"73",
						   57300 => x"F6",		-- 00dfd4: F623             JNE     (mpyl_add_loop)
						   57301 => x"03",
						   57302 => x"0C",		-- 00dfd6: 0C93             TST.W   R12
						   57303 => x"73",
						   57304 => x"F4",		-- 00dfd8: F423             JNE     (mpyl_add_loop)
						   57305 => x"03",
						   57306 => x"0C",		-- 00dfda: 0C4A             MOV.W   R10,R12
						   57307 => x"2A",
						   57308 => x"0D",		-- 00dfdc: 0D4B             MOV.W   R11,R13
						   57309 => x"2B",
						   57310 => x"3A",		-- 00dfde: 3A41             POP.W   R10
						   57311 => x"21",
						   57312 => x"30",		-- 00dfe0: 3041             RET     
						   57313 => x"21",
						   -- Begin: write
						   57314 => x"0C",		-- 00dfe2: 0C93             TST.W   R12
						   57315 => x"73",
						   57316 => x"0E",		-- 00dfe4: 0E38             JL      ($C$L1)
						   57317 => x"18",
						   57318 => x"3C",		-- 00dfe6: 3C90             CMP.W   #0x000a,R12
						   57319 => x"70",
						   57320 => x"0A",		-- 00dfe8: 0A00            
						   57321 => x"00",
						   57322 => x"0B",		-- 00dfea: 0B34             JGE     ($C$L1)
						   57323 => x"14",
						   57324 => x"0C",		-- 00dfec: 0C5C             RLA.W   R12
						   57325 => x"3C",
						   57326 => x"0C",		-- 00dfee: 0C5C             RLA.W   R12
						   57327 => x"3C",
						   57328 => x"3C",		-- 00dff0: 3C50             ADD.W   #0x20c6,R12
						   57329 => x"30",
						   57330 => x"C6",		-- 00dff2: C620            
						   57331 => x"20",
						   57332 => x"2F",		-- 00dff4: 2F4C             MOV.W   @R12,R15
						   57333 => x"2C",
						   57334 => x"0F",		-- 00dff6: 0F93             TST.W   R15
						   57335 => x"73",
						   57336 => x"04",		-- 00dff8: 0424             JEQ     ($C$L1)
						   57337 => x"04",
						   57338 => x"1C",		-- 00dffa: 1C4C             MOV.W   0x0002(R12),R12
						   57339 => x"2C",
						   57340 => x"02",		-- 00dffc: 0200            
						   57341 => x"00",
						   57342 => x"10",		-- 00dffe: 104F             BR      0x0012(R15)
						   57343 => x"2F",
						   57344 => x"12",		-- 00e000: 1200            
						   57345 => x"00",
						   57346 => x"3C",		-- 00e002: 3C43             MOV.W   #-1,R12
						   57347 => x"23",
						   57348 => x"30",		-- 00e004: 3041             RET     
						   57349 => x"21",
						   -- Begin: __mspabi_mpyul
						   -- Begin: __mspabi_mpyul_sw
						   57350 => x"0B",		-- 00e006: 0B4C             MOV.W   R12,R11
						   57351 => x"2C",
						   57352 => x"0E",		-- 00e008: 0E4D             MOV.W   R13,R14
						   57353 => x"2D",
						   57354 => x"0F",		-- 00e00a: 0F43             CLR.W   R15
						   57355 => x"23",
						   57356 => x"0C",		-- 00e00c: 0C43             CLR.W   R12
						   57357 => x"23",
						   57358 => x"0D",		-- 00e00e: 0D43             CLR.W   R13
						   57359 => x"23",
						   57360 => x"12",		-- 00e010: 12C3             CLRC    
						   57361 => x"A3",
						   57362 => x"0B",		-- 00e012: 0B10             RRC     R11
						   57363 => x"F0",
						   57364 => x"01",		-- 00e014: 013C             JMP     (mpyul_add_loop1)
						   57365 => x"1C",
						   -- Begin: mpyul_add_loop
						   57366 => x"0B",		-- 00e016: 0B11             RRA     R11
						   57367 => x"F1",
						   -- Begin: mpyul_add_loop1
						   57368 => x"02",		-- 00e018: 0228             JLO     (shift_test_mpyul)
						   57369 => x"08",
						   57370 => x"0C",		-- 00e01a: 0C5E             ADD.W   R14,R12
						   57371 => x"3E",
						   57372 => x"0D",		-- 00e01c: 0D6F             ADDC.W  R15,R13
						   57373 => x"4F",
						   -- Begin: shift_test_mpyul
						   57374 => x"0E",		-- 00e01e: 0E5E             RLA.W   R14
						   57375 => x"3E",
						   57376 => x"0F",		-- 00e020: 0F6F             RLC.W   R15
						   57377 => x"4F",
						   57378 => x"0B",		-- 00e022: 0B93             TST.W   R11
						   57379 => x"73",
						   57380 => x"F8",		-- 00e024: F823             JNE     (mpyul_add_loop)
						   57381 => x"03",
						   57382 => x"30",		-- 00e026: 3041             RET     
						   57383 => x"21",
						   -- Begin: memccpy
						   57384 => x"0A",		-- 00e028: 0A12             PUSH    R10
						   57385 => x"F2",
						   57386 => x"0F",		-- 00e02a: 0F93             TST.W   R15
						   57387 => x"73",
						   57388 => x"0B",		-- 00e02c: 0B24             JEQ     ($C$L2)
						   57389 => x"04",
						   57390 => x"4E",		-- 00e02e: 4E4E             MOV.B   R14,R14
						   57391 => x"2E",
						   57392 => x"6B",		-- 00e030: 6B4D             MOV.B   @R13,R11
						   57393 => x"2D",
						   57394 => x"1C",		-- 00e032: 1C53             INC.W   R12
						   57395 => x"33",
						   57396 => x"CC",		-- 00e034: CC4B             MOV.B   R11,0xffff(R12)
						   57397 => x"2B",
						   57398 => x"FF",		-- 00e036: FFFF            
						   57399 => x"FF",
						   57400 => x"4A",		-- 00e038: 4A4E             MOV.B   R14,R10
						   57401 => x"2E",
						   57402 => x"0B",		-- 00e03a: 0B9A             CMP.W   R10,R11
						   57403 => x"7A",
						   57404 => x"04",		-- 00e03c: 0424             JEQ     ($C$L3)
						   57405 => x"04",
						   57406 => x"1D",		-- 00e03e: 1D53             INC.W   R13
						   57407 => x"33",
						   57408 => x"1F",		-- 00e040: 1F83             DEC.W   R15
						   57409 => x"63",
						   57410 => x"F6",		-- 00e042: F623             JNE     ($C$L1)
						   57411 => x"03",
						   57412 => x"0C",		-- 00e044: 0C43             CLR.W   R12
						   57413 => x"23",
						   57414 => x"3A",		-- 00e046: 3A41             POP.W   R10
						   57415 => x"21",
						   57416 => x"30",		-- 00e048: 3041             RET     
						   57417 => x"21",
						   -- Begin: __mspabi_mpyull
						   -- Begin: __mspabi_mpyull_sw
						   57418 => x"0A",		-- 00e04a: 0A12             PUSH    R10
						   57419 => x"F2",
						   57420 => x"09",		-- 00e04c: 0912             PUSH    R9
						   57421 => x"F2",
						   57422 => x"08",		-- 00e04e: 0812             PUSH    R8
						   57423 => x"F2",
						   57424 => x"08",		-- 00e050: 084C             MOV.W   R12,R8
						   57425 => x"2C",
						   57426 => x"09",		-- 00e052: 094D             MOV.W   R13,R9
						   57427 => x"2D",
						   57428 => x"0A",		-- 00e054: 0A43             CLR.W   R10
						   57429 => x"23",
						   57430 => x"0B",		-- 00e056: 0B43             CLR.W   R11
						   57431 => x"23",
						   57432 => x"0C",		-- 00e058: 0C4E             MOV.W   R14,R12
						   57433 => x"2E",
						   57434 => x"0D",		-- 00e05a: 0D4F             MOV.W   R15,R13
						   57435 => x"2F",
						   57436 => x"0E",		-- 00e05c: 0E43             CLR.W   R14
						   57437 => x"23",
						   57438 => x"0F",		-- 00e05e: 0F43             CLR.W   R15
						   57439 => x"23",
						   57440 => x"B0",		-- 00e060: B012             CALL    #__mspabi_mpyll_sw
						   57441 => x"F2",
						   57442 => x"EE",		-- 00e062: EEC5            
						   57443 => x"C5",
						   57444 => x"30",		-- 00e064: 3040             BR      #__mspabi_func_epilog_3
						   57445 => x"20",
						   57446 => x"9C",		-- 00e066: 9CE1            
						   57447 => x"E1",
						   -- Begin: _c_int00_noargs
						   57448 => x"31",		-- 00e068: 3140             MOV.W   #0x3000,SP
						   57449 => x"20",
						   57450 => x"00",		-- 00e06a: 0030            
						   57451 => x"30",
						   57452 => x"B0",		-- 00e06c: B012             CALL    #_system_pre_init
						   57453 => x"F2",
						   57454 => x"FC",		-- 00e06e: FCE1            
						   57455 => x"E1",
						   57456 => x"0C",		-- 00e070: 0C93             TST.W   R12
						   57457 => x"73",
						   57458 => x"02",		-- 00e072: 0224             JEQ     ($C$L2)
						   57459 => x"04",
						   57460 => x"B0",		-- 00e074: B012             CALL    #__TI_auto_init_nobinit_nopinit
						   57461 => x"F2",
						   57462 => x"D8",		-- 00e076: D8DB            
						   57463 => x"DB",
						   57464 => x"0C",		-- 00e078: 0C43             CLR.W   R12
						   57465 => x"23",
						   57466 => x"B0",		-- 00e07a: B012             CALL    #main
						   57467 => x"F2",
						   57468 => x"3C",		-- 00e07c: 3CD8            
						   57469 => x"D8",
						   57470 => x"1C",		-- 00e07e: 1C43             MOV.W   #1,R12
						   57471 => x"23",
						   57472 => x"B0",		-- 00e080: B012             CALL    #exit
						   57473 => x"F2",
						   57474 => x"94",		-- 00e082: 94DB            
						   57475 => x"DB",
						   -- Begin: free_list_remove
						   57476 => x"3F",		-- 00e084: 3F40             MOV.W   #0x21a6,R15
						   57477 => x"20",
						   57478 => x"A6",		-- 00e086: A621            
						   57479 => x"21",
						   57480 => x"02",		-- 00e088: 023C             JMP     ($C$L2)
						   57481 => x"1C",
						   57482 => x"2F",		-- 00e08a: 2F42             MOV.W   #4,R15
						   57483 => x"22",
						   57484 => x"0F",		-- 00e08c: 0F5E             ADD.W   R14,R15
						   57485 => x"3E",
						   57486 => x"2E",		-- 00e08e: 2E4F             MOV.W   @R15,R14
						   57487 => x"2F",
						   57488 => x"0E",		-- 00e090: 0E93             TST.W   R14
						   57489 => x"73",
						   57490 => x"05",		-- 00e092: 0524             JEQ     ($C$L3)
						   57491 => x"04",
						   57492 => x"0E",		-- 00e094: 0E9C             CMP.W   R12,R14
						   57493 => x"7C",
						   57494 => x"F9",		-- 00e096: F923             JNE     ($C$L1)
						   57495 => x"03",
						   57496 => x"9F",		-- 00e098: 9F4C             MOV.W   0x0004(R12),0x0000(R15)
						   57497 => x"2C",
						   57498 => x"04",		-- 00e09a: 0400            
						   57499 => x"00",
						   57500 => x"00",		-- 00e09c: 0000            
						   57501 => x"00",
						   57502 => x"30",		-- 00e09e: 3041             RET     
						   57503 => x"21",
						   -- Begin: strchr
						   57504 => x"6F",		-- 00e0a0: 6F4C             MOV.B   @R12,R15
						   57505 => x"2C",
						   57506 => x"4D",		-- 00e0a2: 4D4D             MOV.B   R13,R13
						   57507 => x"2D",
						   57508 => x"06",		-- 00e0a4: 063C             JMP     ($C$L3)
						   57509 => x"1C",
						   57510 => x"0F",		-- 00e0a6: 0F93             TST.W   R15
						   57511 => x"73",
						   57512 => x"02",		-- 00e0a8: 0220             JNE     ($C$L2)
						   57513 => x"00",
						   57514 => x"0C",		-- 00e0aa: 0C43             CLR.W   R12
						   57515 => x"23",
						   57516 => x"30",		-- 00e0ac: 3041             RET     
						   57517 => x"21",
						   57518 => x"1C",		-- 00e0ae: 1C53             INC.W   R12
						   57519 => x"33",
						   57520 => x"6F",		-- 00e0b0: 6F4C             MOV.B   @R12,R15
						   57521 => x"2C",
						   57522 => x"4E",		-- 00e0b2: 4E4D             MOV.B   R13,R14
						   57523 => x"2D",
						   57524 => x"0F",		-- 00e0b4: 0F9E             CMP.W   R14,R15
						   57525 => x"7E",
						   57526 => x"F7",		-- 00e0b6: F723             JNE     ($C$L1)
						   57527 => x"03",
						   57528 => x"30",		-- 00e0b8: 3041             RET     
						   57529 => x"21",
						   -- Begin: strcmp
						   57530 => x"0F",		-- 00e0ba: 0F4C             MOV.W   R12,R15
						   57531 => x"2C",
						   57532 => x"6E",		-- 00e0bc: 6E4F             MOV.B   @R15,R14
						   57533 => x"2F",
						   57534 => x"6B",		-- 00e0be: 6B4D             MOV.B   @R13,R11
						   57535 => x"2D",
						   57536 => x"4C",		-- 00e0c0: 4C4E             MOV.B   R14,R12
						   57537 => x"2E",
						   57538 => x"0C",		-- 00e0c2: 0C8B             SUB.W   R11,R12
						   57539 => x"6B",
						   57540 => x"4E",		-- 00e0c4: 4E93             TST.B   R14
						   57541 => x"73",
						   57542 => x"04",		-- 00e0c6: 0424             JEQ     ($C$L2)
						   57543 => x"04",
						   57544 => x"1D",		-- 00e0c8: 1D53             INC.W   R13
						   57545 => x"33",
						   57546 => x"1F",		-- 00e0ca: 1F53             INC.W   R15
						   57547 => x"33",
						   57548 => x"0C",		-- 00e0cc: 0C93             TST.W   R12
						   57549 => x"73",
						   57550 => x"F6",		-- 00e0ce: F627             JEQ     ($C$L1)
						   57551 => x"07",
						   57552 => x"30",		-- 00e0d0: 3041             RET     
						   57553 => x"21",
						   -- Begin: __mspabi_divu
						   -- Begin: __mspabi_remu
						   57554 => x"0E",		-- 00e0d2: 0E43             CLR.W   R14
						   57555 => x"23",
						   57556 => x"0F",		-- 00e0d4: 0F4C             MOV.W   R12,R15
						   57557 => x"2C",
						   57558 => x"1C",		-- 00e0d6: 1C43             MOV.W   #1,R12
						   57559 => x"23",
						   -- Begin: div_loop
						   57560 => x"0F",		-- 00e0d8: 0F5F             RLA.W   R15
						   57561 => x"3F",
						   57562 => x"0E",		-- 00e0da: 0E6E             RLC.W   R14
						   57563 => x"4E",
						   57564 => x"0E",		-- 00e0dc: 0E9D             CMP.W   R13,R14
						   57565 => x"7D",
						   57566 => x"01",		-- 00e0de: 0128             JLO     (set_quotient_bit)
						   57567 => x"08",
						   57568 => x"0E",		-- 00e0e0: 0E8D             SUB.W   R13,R14
						   57569 => x"6D",
						   -- Begin: set_quotient_bit
						   57570 => x"0C",		-- 00e0e2: 0C6C             RLC.W   R12
						   57571 => x"4C",
						   57572 => x"F9",		-- 00e0e4: F92B             JLO     (div_loop)
						   57573 => x"0B",
						   57574 => x"30",		-- 00e0e6: 3041             RET     
						   57575 => x"21",
						   -- Begin: __TI_zero_init_nomemset
						   57576 => x"1F",		-- 00e0e8: 1F4C             MOV.W   0x0001(R12),R15
						   57577 => x"2C",
						   57578 => x"01",		-- 00e0ea: 0100            
						   57579 => x"00",
						   57580 => x"0F",		-- 00e0ec: 0F93             TST.W   R15
						   57581 => x"73",
						   57582 => x"05",		-- 00e0ee: 0524             JEQ     ($C$L2)
						   57583 => x"04",
						   57584 => x"1D",		-- 00e0f0: 1D53             INC.W   R13
						   57585 => x"33",
						   57586 => x"CD",		-- 00e0f2: CD43             CLR.B   0xffff(R13)
						   57587 => x"23",
						   57588 => x"FF",		-- 00e0f4: FFFF            
						   57589 => x"FF",
						   57590 => x"1F",		-- 00e0f6: 1F83             DEC.W   R15
						   57591 => x"63",
						   57592 => x"FB",		-- 00e0f8: FB23             JNE     ($C$L1)
						   57593 => x"03",
						   57594 => x"30",		-- 00e0fa: 3041             RET     
						   57595 => x"21",
						   -- Begin: memchr
						   57596 => x"0E",		-- 00e0fc: 0E93             TST.W   R14
						   57597 => x"73",
						   57598 => x"06",		-- 00e0fe: 0624             JEQ     ($C$L2)
						   57599 => x"04",
						   57600 => x"4D",		-- 00e100: 4D4D             MOV.B   R13,R13
						   57601 => x"2D",
						   57602 => x"6D",		-- 00e102: 6D9C             CMP.B   @R12,R13
						   57603 => x"7C",
						   57604 => x"04",		-- 00e104: 0424             JEQ     ($C$L3)
						   57605 => x"04",
						   57606 => x"1C",		-- 00e106: 1C53             INC.W   R12
						   57607 => x"33",
						   57608 => x"1E",		-- 00e108: 1E83             DEC.W   R14
						   57609 => x"63",
						   57610 => x"FB",		-- 00e10a: FB23             JNE     ($C$L1)
						   57611 => x"03",
						   57612 => x"0C",		-- 00e10c: 0C43             CLR.W   R12
						   57613 => x"23",
						   57614 => x"30",		-- 00e10e: 3041             RET     
						   57615 => x"21",
						   -- Begin: memset
						   57616 => x"0F",		-- 00e110: 0F4C             MOV.W   R12,R15
						   57617 => x"2C",
						   57618 => x"0E",		-- 00e112: 0E93             TST.W   R14
						   57619 => x"73",
						   57620 => x"06",		-- 00e114: 0624             JEQ     ($C$L2)
						   57621 => x"04",
						   57622 => x"4D",		-- 00e116: 4D4D             MOV.B   R13,R13
						   57623 => x"2D",
						   57624 => x"1F",		-- 00e118: 1F53             INC.W   R15
						   57625 => x"33",
						   57626 => x"CF",		-- 00e11a: CF4D             MOV.B   R13,0xffff(R15)
						   57627 => x"2D",
						   57628 => x"FF",		-- 00e11c: FFFF            
						   57629 => x"FF",
						   57630 => x"1E",		-- 00e11e: 1E83             DEC.W   R14
						   57631 => x"63",
						   57632 => x"FB",		-- 00e120: FB23             JNE     ($C$L1)
						   57633 => x"03",
						   57634 => x"30",		-- 00e122: 3041             RET     
						   57635 => x"21",
						   -- Begin: __mspabi_mpyi
						   -- Begin: __mspabi_mpyi_sw
						   57636 => x"0E",		-- 00e124: 0E43             CLR.W   R14
						   57637 => x"23",
						   -- Begin: mpyi_add_loop
						   57638 => x"12",		-- 00e126: 12C3             CLRC    
						   57639 => x"A3",
						   57640 => x"0C",		-- 00e128: 0C10             RRC     R12
						   57641 => x"F0",
						   57642 => x"01",		-- 00e12a: 0128             JLO     (shift_test_mpyi)
						   57643 => x"08",
						   57644 => x"0E",		-- 00e12c: 0E5D             ADD.W   R13,R14
						   57645 => x"3D",
						   -- Begin: shift_test_mpyi
						   57646 => x"0D",		-- 00e12e: 0D5D             RLA.W   R13
						   57647 => x"3D",
						   57648 => x"0C",		-- 00e130: 0C93             TST.W   R12
						   57649 => x"73",
						   57650 => x"F9",		-- 00e132: F923             JNE     (mpyi_add_loop)
						   57651 => x"03",
						   57652 => x"0C",		-- 00e134: 0C4E             MOV.W   R14,R12
						   57653 => x"2E",
						   57654 => x"30",		-- 00e136: 3041             RET     
						   57655 => x"21",
						   -- Begin: wcslen
						   57656 => x"0F",		-- 00e138: 0F4C             MOV.W   R12,R15
						   57657 => x"2C",
						   57658 => x"01",		-- 00e13a: 013C             JMP     ($C$L2)
						   57659 => x"1C",
						   57660 => x"2F",		-- 00e13c: 2F53             INCD.W  R15
						   57661 => x"33",
						   57662 => x"8F",		-- 00e13e: 8F93             TST.W   0x0000(R15)
						   57663 => x"73",
						   57664 => x"00",		-- 00e140: 0000            
						   57665 => x"00",
						   57666 => x"FC",		-- 00e142: FC23             JNE     ($C$L1)
						   57667 => x"03",
						   57668 => x"0F",		-- 00e144: 0F8C             SUB.W   R12,R15
						   57669 => x"6C",
						   57670 => x"0F",		-- 00e146: 0F11             RRA     R15
						   57671 => x"F1",
						   57672 => x"0C",		-- 00e148: 0C4F             MOV.W   R15,R12
						   57673 => x"2F",
						   57674 => x"30",		-- 00e14a: 3041             RET     
						   57675 => x"21",
						   -- Begin: buff_value
						   57676 => x"21",		-- 00e14c: 2183             DECD.W  SP
						   57677 => x"63",
						   57678 => x"81",		-- 00e14e: 814C             MOV.W   R12,0x0000(SP)
						   57679 => x"2C",
						   57680 => x"00",		-- 00e150: 0000            
						   57681 => x"00",
						   57682 => x"3D",		-- 00e152: 3D40             MOV.W   #0x8514,R13
						   57683 => x"20",
						   57684 => x"14",		-- 00e154: 1485            
						   57685 => x"85",
						   57686 => x"B0",		-- 00e156: B012             CALL    #strcpy
						   57687 => x"F2",
						   57688 => x"A4",		-- 00e158: A4E1            
						   57689 => x"E1",
						   57690 => x"21",		-- 00e15a: 2153             INCD.W  SP
						   57691 => x"33",
						   57692 => x"30",		-- 00e15c: 3041             RET     
						   57693 => x"21",
						   -- Begin: __TI_decompress_none
						   57694 => x"0F",		-- 00e15e: 0F4C             MOV.W   R12,R15
						   57695 => x"2C",
						   57696 => x"0C",		-- 00e160: 0C4D             MOV.W   R13,R12
						   57697 => x"2D",
						   57698 => x"3D",		-- 00e162: 3D40             MOV.W   #0x0003,R13
						   57699 => x"20",
						   57700 => x"03",		-- 00e164: 0300            
						   57701 => x"00",
						   57702 => x"0D",		-- 00e166: 0D5F             ADD.W   R15,R13
						   57703 => x"3F",
						   57704 => x"1E",		-- 00e168: 1E4F             MOV.W   0x0001(R15),R14
						   57705 => x"2F",
						   57706 => x"01",		-- 00e16a: 0100            
						   57707 => x"00",
						   57708 => x"30",		-- 00e16c: 3040             BR      #memcpy
						   57709 => x"20",
						   57710 => x"82",		-- 00e16e: 82E1            
						   57711 => x"E1",
						   -- Begin: __mspabi_srll
						   57712 => x"3E",		-- 00e170: 3EF0             AND.W   #0x001f,R14
						   57713 => x"D0",
						   57714 => x"1F",		-- 00e172: 1F00            
						   57715 => x"00",
						   57716 => x"05",		-- 00e174: 0524             JEQ     (L_LSR_RET)
						   57717 => x"04",
						   -- Begin: L_LSR_TOP
						   57718 => x"12",		-- 00e176: 12C3             CLRC    
						   57719 => x"A3",
						   57720 => x"0D",		-- 00e178: 0D10             RRC     R13
						   57721 => x"F0",
						   57722 => x"0C",		-- 00e17a: 0C10             RRC     R12
						   57723 => x"F0",
						   57724 => x"1E",		-- 00e17c: 1E83             DEC.W   R14
						   57725 => x"63",
						   57726 => x"FB",		-- 00e17e: FB23             JNE     (L_LSR_TOP)
						   57727 => x"03",
						   -- Begin: L_LSR_RET
						   57728 => x"30",		-- 00e180: 3041             RET     
						   57729 => x"21",
						   -- Begin: memcpy
						   57730 => x"0E",		-- 00e182: 0E93             TST.W   R14
						   57731 => x"73",
						   57732 => x"06",		-- 00e184: 0624             JEQ     ($C$L2)
						   57733 => x"04",
						   57734 => x"0F",		-- 00e186: 0F4C             MOV.W   R12,R15
						   57735 => x"2C",
						   57736 => x"1F",		-- 00e188: 1F53             INC.W   R15
						   57737 => x"33",
						   57738 => x"FF",		-- 00e18a: FF4D             MOV.B   @R13+,0xffff(R15)
						   57739 => x"2D",
						   57740 => x"FF",		-- 00e18c: FFFF            
						   57741 => x"FF",
						   57742 => x"1E",		-- 00e18e: 1E83             DEC.W   R14
						   57743 => x"63",
						   57744 => x"FB",		-- 00e190: FB23             JNE     ($C$L1)
						   57745 => x"03",
						   57746 => x"30",		-- 00e192: 3041             RET     
						   57747 => x"21",
						   -- Begin: __mspabi_func_epilog_7
						   -- Begin: __mspabi_func_epilog
						   57748 => x"34",		-- 00e194: 3441             POP.W   R4
						   57749 => x"21",
						   -- Begin: __mspabi_func_epilog_6
						   57750 => x"35",		-- 00e196: 3541             POP.W   R5
						   57751 => x"21",
						   -- Begin: __mspabi_func_epilog_5
						   57752 => x"36",		-- 00e198: 3641             POP.W   R6
						   57753 => x"21",
						   -- Begin: __mspabi_func_epilog_4
						   57754 => x"37",		-- 00e19a: 3741             POP.W   R7
						   57755 => x"21",
						   -- Begin: __mspabi_func_epilog_3
						   57756 => x"38",		-- 00e19c: 3841             POP.W   R8
						   57757 => x"21",
						   -- Begin: __mspabi_func_epilog_2
						   57758 => x"39",		-- 00e19e: 3941             POP.W   R9
						   57759 => x"21",
						   -- Begin: __mspabi_func_epilog_1
						   57760 => x"3A",		-- 00e1a0: 3A41             POP.W   R10
						   57761 => x"21",
						   57762 => x"30",		-- 00e1a2: 3041             RET     
						   57763 => x"21",
						   -- Begin: strcpy
						   57764 => x"0F",		-- 00e1a4: 0F4C             MOV.W   R12,R15
						   57765 => x"2C",
						   57766 => x"7E",		-- 00e1a6: 7E4D             MOV.B   @R13+,R14
						   57767 => x"2D",
						   57768 => x"1F",		-- 00e1a8: 1F53             INC.W   R15
						   57769 => x"33",
						   57770 => x"CF",		-- 00e1aa: CF4E             MOV.B   R14,0xffff(R15)
						   57771 => x"2E",
						   57772 => x"FF",		-- 00e1ac: FFFF            
						   57773 => x"FF",
						   57774 => x"0E",		-- 00e1ae: 0E93             TST.W   R14
						   57775 => x"73",
						   57776 => x"FA",		-- 00e1b0: FA23             JNE     ($C$L1)
						   57777 => x"03",
						   57778 => x"30",		-- 00e1b2: 3041             RET     
						   57779 => x"21",
						   -- Begin: strlen
						   57780 => x"3F",		-- 00e1b4: 3F43             MOV.W   #-1,R15
						   57781 => x"23",
						   57782 => x"1F",		-- 00e1b6: 1F53             INC.W   R15
						   57783 => x"33",
						   57784 => x"7E",		-- 00e1b8: 7E4C             MOV.B   @R12+,R14
						   57785 => x"2C",
						   57786 => x"0E",		-- 00e1ba: 0E93             TST.W   R14
						   57787 => x"73",
						   57788 => x"FC",		-- 00e1bc: FC23             JNE     ($C$L1)
						   57789 => x"03",
						   57790 => x"0C",		-- 00e1be: 0C4F             MOV.W   R15,R12
						   57791 => x"2F",
						   57792 => x"30",		-- 00e1c0: 3041             RET     
						   57793 => x"21",
						   -- Begin: __mspabi_fltid
						   57794 => x"3C",		-- 00e1c2: 3CB0             BIT.W   #0x8000,R12
						   57795 => x"90",
						   57796 => x"00",		-- 00e1c4: 0080            
						   57797 => x"80",
						   57798 => x"0D",		-- 00e1c6: 0D7D             SUBC.W  R13,R13
						   57799 => x"5D",
						   57800 => x"3D",		-- 00e1c8: 3DE3             INV.W   R13
						   57801 => x"C3",
						   57802 => x"30",		-- 00e1ca: 3040             BR      #__mspabi_fltlid
						   57803 => x"20",
						   57804 => x"AC",		-- 00e1cc: ACCE            
						   57805 => x"CE",
						   -- Begin: toupper
						   57806 => x"EC",		-- 00e1ce: ECB3             BIT.B   #2,0x992f(R12)
						   57807 => x"93",
						   57808 => x"2F",		-- 00e1d0: 2F99            
						   57809 => x"99",
						   57810 => x"02",		-- 00e1d2: 0224             JEQ     ($C$L1)
						   57811 => x"04",
						   57812 => x"3C",		-- 00e1d4: 3C80             SUB.W   #0x0020,R12
						   57813 => x"60",
						   57814 => x"20",		-- 00e1d6: 2000            
						   57815 => x"00",
						   57816 => x"30",		-- 00e1d8: 3041             RET     
						   57817 => x"21",
						   -- Begin: abs
						   57818 => x"0C",		-- 00e1da: 0C93             TST.W   R12
						   57819 => x"73",
						   57820 => x"02",		-- 00e1dc: 0234             JGE     ($C$L1)
						   57821 => x"14",
						   57822 => x"3C",		-- 00e1de: 3CE3             INV.W   R12
						   57823 => x"C3",
						   57824 => x"1C",		-- 00e1e0: 1C53             INC.W   R12
						   57825 => x"33",
						   57826 => x"30",		-- 00e1e2: 3041             RET     
						   57827 => x"21",
						   -- Begin: malloc
						   57828 => x"0D",		-- 00e1e4: 0D4C             MOV.W   R12,R13
						   57829 => x"2C",
						   57830 => x"2C",		-- 00e1e6: 2C42             MOV.W   #4,R12
						   57831 => x"22",
						   57832 => x"30",		-- 00e1e8: 3040             BR      #aligned_alloc
						   57833 => x"20",
						   57834 => x"FA",		-- 00e1ea: FAC7            
						   57835 => x"C7",
						   -- Begin: _outc
						   57836 => x"4C",		-- 00e1ec: 4C4C             MOV.B   R12,R12
						   57837 => x"2C",
						   57838 => x"30",		-- 00e1ee: 3040             BR      #fputc
						   57839 => x"20",
						   57840 => x"96",		-- 00e1f0: 96D0            
						   57841 => x"D0",
						   -- Begin: abort
						   57842 => x"03",		-- 00e1f2: 0343             NOP     
						   57843 => x"23",
						   57844 => x"FF",		-- 00e1f4: FF3F             JMP     ($C$L1)
						   57845 => x"1F",
						   57846 => x"03",		-- 00e1f6: 0343             NOP     
						   57847 => x"23",
						   -- Begin: _outs
						   57848 => x"30",		-- 00e1f8: 3040             BR      #fputs
						   57849 => x"20",
						   57850 => x"F0",		-- 00e1fa: F0C8            
						   57851 => x"C8",
						   -- Begin: _system_pre_init
						   57852 => x"1C",		-- 00e1fc: 1C43             MOV.W   #1,R12
						   57853 => x"23",
						   57854 => x"30",		-- 00e1fe: 3041             RET     
						   57855 => x"21",
						   -- Begin: _nop
						   57856 => x"30",		-- 00e200: 3041             RET     
						   57857 => x"21",
						   -- Begin: _system_post_cinit
						   57858 => x"30",		-- 00e202: 3041             RET     
						   57859 => x"21",
						   -- ISR Trap
						   57860 => x"32",		-- 00e204: 32D0             BIS.W   #0x0010,SR
						   57861 => x"B0",
						   57862 => x"10",		-- 00e206: 1000            
						   57863 => x"00",
						   57864 => x"FD",		-- 00e208: FD3F             JMP     (__TI_ISR_TRAP)
						   57865 => x"1F",
						   57866 => x"03",		-- 00e20a: 0343             NOP     
						   57867 => x"23",
						   -- IRQ Vectors (Interrupt Vectors)
						   65486 => x"04",		-- 00ffce:e204 PORT4 __TI_int22 int22
						   65487 => x"e2",
						   65488 => x"04",		-- 00ffd0:e204 PORT3 __TI_int23 int23
						   65489 => x"e2",
						   65490 => x"04",		-- 00ffd2:e204 PORT2 __TI_int24 int24
						   65491 => x"e2",
						   65492 => x"04",		-- 00ffd4:e204 PORT1 __TI_int25 int25
						   65493 => x"e2",
						   65494 => x"04",		-- 00ffd6:e204 SAC1_SAC3 __TI_int26 int26
						   65495 => x"e2",
						   65496 => x"04",		-- 00ffd8:e204 SAC0_SAC2 __TI_int27 int27
						   65497 => x"e2",
						   65498 => x"04",		-- 00ffda:e204 ECOMP0_ECOMP1 __TI_int28 int28
						   65499 => x"e2",
						   65500 => x"04",		-- 00ffdc:e204 ADC __TI_int29 int29
						   65501 => x"e2",
						   65502 => x"04",		-- 00ffde:e204 EUSCI_B1 __TI_int30 int30
						   65503 => x"e2",
						   65504 => x"04",		-- 00ffe0:e204 EUSCI_B0 __TI_int31 int31
						   65505 => x"e2",
						   65506 => x"04",		-- 00ffe2:e204 EUSCI_A1 __TI_int32 int32
						   65507 => x"e2",
						   65508 => x"04",		-- 00ffe4:e204 EUSCI_A0 __TI_int33 int33
						   65509 => x"e2",
						   65510 => x"04",		-- 00ffe6:e204 WDT __TI_int34 int34
						   65511 => x"e2",
						   65512 => x"04",		-- 00ffe8:e204 RTC __TI_int35 int35
						   65513 => x"e2",
						   65514 => x"04",		-- 00ffea:e204 TIMER3_B1 __TI_int36 int36
						   65515 => x"e2",
						   65516 => x"04",		-- 00ffec:e204 TIMER3_B0 __TI_int37 int37
						   65517 => x"e2",
						   65518 => x"04",		-- 00ffee:e204 TIMER2_B1 __TI_int38 int38
						   65519 => x"e2",
						   65520 => x"04",		-- 00fff0:e204 TIMER2_B0 __TI_int39 int39
						   65521 => x"e2",
						   65522 => x"04",		-- 00fff2:e204 TIMER1_B1 __TI_int40 int40
						   65523 => x"e2",
						   65524 => x"04",		-- 00fff4:e204 TIMER1_B0 __TI_int41 int41
						   65525 => x"e2",
						   65526 => x"04",		-- 00fff6:e204 TIMER0_B1 __TI_int42 int42
						   65527 => x"e2",
						   65528 => x"04",		-- 00fff8:e204 TIMER0_B0 __TI_int43 int43
						   65529 => x"e2",
						   65530 => x"04",		-- 00fffa:e204 UNMI __TI_int44 int44
						   65531 => x"e2",
						   65532 => x"04",		-- 00fffc:e204 SYSNMI __TI_int45 int45
						   65533 => x"e2",

                           65534 =>  x"00",		-- Reset Vector = xFFFE:xFFFF
                           65535 =>  x"80",		--  Startup Value = x8000

                           others => x"00");

    signal EN : std_logic;
    
    begin
    -- Note 1:  The bus system uses a 16-bit Address (MAB)
    --          This address size can access locations from x0000 to xFFFF
    --          But our array is only defined from x8000 to xFFFF and
    --          if we try to access it with any other address, it will crash.
    --          So the first thing we need to do is create a local enable that
    --          will only assert when MAB is within x8000 to xFFFF.

     LOCAL_EN : process (MAB) 
     begin
         if ( (to_integer(unsigned(MAB)) >= 32768) and (to_integer(unsigned(MAB)) <= 65535)) then
           EN <= '1';
         else 
           EN <= '0';
         end if;
     end process;

    
    -- Note 2:  The bus system uses a 16-bit Address (MAB)
    --          The MDB_out is also provided as a 16-bit word
    --          However, the memory array is actually built as 8-bit bytes.
    --          So for a given 16-bit MAB, we give MDB_out = HB : LB
    --                                                 or  = ROM(MAB);1) : ROM(MAB)

    MEMORY_ROM : process (clk) 
    begin
        if (rising_edge(clk)) then
            if (EN='1' and write='0') then                      
              MDB_in <= ROM(to_integer(unsigned(MAB)) + 1 ) & ROM(to_integer(unsigned(MAB))); 
            end if;
        end if;
    end process;


end architecture;